module pyramid_synthetic_exposure_fusion_opt(
	input clk,
	input rst,
	input start,
	output done,
	logic [0:0] buf_in_off_chip_clk,
	logic [0:0] buf_in_off_chip_rst,
	logic [0:0] buf_in_off_chip_start,
	logic [0:0] buf_in_off_chip_done,
	logic [31:0] buf_in_off_chip_in_update_0_read_dummy,
	logic [0:0] buf_in_off_chip_in_off_chip_update_0_write_wen,
	logic [31:0] buf_in_off_chip_in_off_chip_update_0_write_wdata,
	logic [31:0] buf_in_off_chip_in_update_0_read_rdata,
	logic [0:0] buf_pyramid_synthetic_exposure_fusion_clk,
	logic [0:0] buf_pyramid_synthetic_exposure_fusion_rst,
	logic [0:0] buf_pyramid_synthetic_exposure_fusion_start,
	logic [0:0] buf_pyramid_synthetic_exposure_fusion_done,
	logic [0:0] buf_pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_wen,
	logic [31:0] buf_pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_wdata);

  logic [31:0] in_off_chip_in_update_0_read_read_0;
  logic [31:0] in_update_0;
  logic [31:0] bright_bright_weights_update_0_read_read_4;
  logic [31:0] bright_weights_update_0;
  logic [31:0] bright_weights_bright_weights_update_0_write_write_5;
  logic [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57;
  logic [31:0] dark_dark_weights_update_0_read_read_8;
  logic [31:0] dark_weights_update_0;
  logic [31:0] dark_weights_dark_weights_update_0_write_write_9;
  logic [31:0] dark_weights_normed_gauss_blur_2_update_0;
  logic [31:0] final_merged_2_final_merged_1_update_0_read_read_120;
  logic [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58;
  logic [31:0] fused_level_1_final_merged_1_update_0_read_read_121;
  logic [31:0] final_merged_1_update_0;
  logic [31:0] final_merged_1_final_merged_1_update_0_write_write_122;
  logic [31:0] in_in_update_0_write_write_1;
  logic [31:0] in_bright_update_0_read_read_2;
  logic [31:0] bright_update_0;
  logic [31:0] bright_bright_update_0_write_write_3;
  logic [31:0] in_dark_update_0_read_read_6;
  logic [31:0] dark_update_0;
  logic [31:0] dark_dark_update_0_write_write_7;
  logic [287:0] dark_dark_gauss_blur_1_update_0_read_read_10;
  logic [31:0] dark_gauss_blur_1_update_0;
  logic [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39;
  logic [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11;
  logic [31:0] bright_gauss_blur_1_update_0;
  logic [287:0] bright_bright_gauss_blur_1_update_0_read_read_12;
  logic [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13;
  logic [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40;
  logic [31:0] bright_laplace_us_1_update_0;
  logic [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41;
  logic [31:0] bright_weights_normed_gauss_blur_1_update_0;
  logic [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55;
  logic [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59;
  logic [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56;
  logic [31:0] bright_laplace_us_2_update_0;
  logic [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60;
  logic [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61;
  logic [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102;
  logic [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114;
  logic [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115;
  logic [31:0] fused_level_3_update_0;
  logic [31:0] fused_level_3_fused_level_3_update_0_write_write_116;
  logic [31:0] fused_level_3_final_merged_2_update_0_read_read_117;
  logic [31:0] fused_level_2_final_merged_2_update_0_read_read_118;
  logic [31:0] final_merged_2_update_0;
  logic [31:0] final_merged_2_final_merged_2_update_0_write_write_119;
  logic [31:0] final_merged_1_final_merged_0_update_0_read_read_123;
  logic [31:0] fused_level_0_final_merged_0_update_0_read_read_124;
  logic [31:0] final_merged_0_update_0;
  logic [31:0] final_merged_0_final_merged_0_update_0_write_write_125;
  logic [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16;
  logic [31:0] dark_laplace_us_0_update_0;
  logic [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17;
  logic [31:0] dark_weights_weight_sums_update_0_read_read_22;
  logic [31:0] weight_sums_update_0;
  logic [31:0] bright_weights_weight_sums_update_0_read_read_23;
  logic [31:0] weight_sums_weight_sums_update_0_write_write_24;
  logic [31:0] dark_dark_laplace_diff_0_update_0_read_read_27;
  logic [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28;
  logic [31:0] dark_laplace_diff_0_update_0;
  logic [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29;
  logic [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32;
  logic [31:0] bright_gauss_ds_2_update_0;
  logic [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38;
  logic [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33;
  logic [31:0] bright_gauss_ds_3_update_0;
  logic [31:0] bright_bright_laplace_diff_0_update_0_read_read_42;
  logic [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43;
  logic [31:0] bright_laplace_diff_0_update_0;
  logic [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44;
  logic [31:0] bright_weights_bright_weights_normed_update_0_read_read_48;
  logic [31:0] weight_sums_bright_weights_normed_update_0_read_read_49;
  logic [31:0] bright_weights_normed_update_0;
  logic [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50;
  logic [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53;
  logic [31:0] dark_weights_normed_gauss_ds_1_update_0;
  logic [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65;
  logic [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54;
  logic [31:0] dark_gauss_blur_3_update_0;
  logic [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66;
  logic [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70;
  logic [31:0] bright_weights_normed_gauss_ds_1_update_0;
  logic [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71;
  logic [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87;
  logic [31:0] fused_level_1_update_0;
  logic [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88;
  logic [31:0] fused_level_1_fused_level_1_update_0_write_write_89;
  logic [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94;
  logic [31:0] dark_weights_normed_gauss_ds_3_update_0;
  logic [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98;
  logic [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95;
  logic [31:0] dark_laplace_us_2_update_0;
  logic [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99;
  logic [31:0] final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126;
  logic [31:0] pyramid_synthetic_exposure_fusion_update_0;
  logic [31:0] pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127;
  logic [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14;
  logic [31:0] dark_gauss_ds_1_update_0;
  logic [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15;
  logic [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19;
  logic [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20;
  logic [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18;
  logic [31:0] dark_gauss_blur_2_update_0;
  logic [31:0] bright_gauss_ds_1_update_0;
  logic [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21;
  logic [31:0] weight_sums_dark_weights_normed_update_0_read_read_46;
  logic [31:0] dark_weights_normed_update_0;
  logic [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25;
  logic [31:0] bright_gauss_blur_2_update_0;
  logic [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26;
  logic [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30;
  logic [31:0] bright_laplace_us_0_update_0;
  logic [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31;
  logic [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34;
  logic [31:0] dark_gauss_ds_2_update_0;
  logic [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35;
  logic [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72;
  logic [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36;
  logic [31:0] bright_gauss_blur_3_update_0;
  logic [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37;
  logic [31:0] dark_weights_dark_weights_normed_update_0_read_read_45;
  logic [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47;
  logic [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51;
  logic [31:0] dark_weights_normed_gauss_blur_1_update_0;
  logic [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52;
  logic [31:0] dark_laplace_us_1_update_0;
  logic [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62;
  logic [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67;
  logic [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63;
  logic [31:0] dark_weights_normed_gauss_ds_2_update_0;
  logic [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64;
  logic [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68;
  logic [31:0] bright_laplace_diff_1_update_0;
  logic [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69;
  logic [31:0] dark_weights_normed_gauss_blur_3_update_0;
  logic [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73;
  logic [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74;
  logic [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75;
  logic [31:0] dark_laplace_diff_1_update_0;
  logic [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76;
  logic [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82;
  logic [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77;
  logic [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78;
  logic [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79;
  logic [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80;
  logic [31:0] fused_level_0_update_0;
  logic [31:0] fused_level_0_fused_level_0_update_0_write_write_81;
  logic [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83;
  logic [31:0] bright_laplace_diff_2_update_0;
  logic [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84;
  logic [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90;
  logic [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85;
  logic [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86;
  logic [31:0] bright_weights_normed_gauss_blur_2_update_0;
  logic [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92;
  logic [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91;
  logic [31:0] dark_gauss_ds_3_update_0;
  logic [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93;
  logic [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96;
  logic [31:0] bright_weights_normed_gauss_ds_2_update_0;
  logic [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97;
  logic [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100;
  logic [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101;
  logic [31:0] dark_laplace_diff_2_update_0;
  logic [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103;
  logic [31:0] bright_weights_normed_gauss_blur_3_update_0;
  logic [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104;
  logic [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105;
  logic [31:0] bright_weights_normed_gauss_ds_3_update_0;
  logic [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107;
  logic [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106;
  logic [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108;
  logic [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109;
  logic [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110;
  logic [31:0] fused_level_2_update_0;
  logic [31:0] fused_level_2_fused_level_2_update_0_write_write_111;
  logic [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112;
  logic [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113;

  logic started;

  logic stage_0_active;
  logic stage_1_active;
  logic stage_2_active;
  logic stage_3_active;
  logic stage_4_active;
  logic stage_5_active;
  logic stage_6_active;
  logic stage_7_active;
  logic stage_8_active;
  logic stage_9_active;
  logic stage_10_active;
  logic stage_11_active;
  logic stage_12_active;
  logic stage_13_active;
  logic stage_14_active;
  logic stage_15_active;
  logic stage_16_active;
  logic stage_17_active;
  logic stage_18_active;
  logic stage_19_active;
  logic stage_20_active;
  logic stage_21_active;
  logic stage_22_active;
  logic stage_23_active;
  logic stage_24_active;
  logic stage_25_active;
  logic stage_26_active;
  logic stage_27_active;
  logic stage_28_active;
  logic stage_29_active;
  logic stage_30_active;
  logic stage_31_active;
  logic stage_32_active;
  logic stage_33_active;
  logic stage_34_active;
  logic stage_35_active;
  logic stage_36_active;
  logic stage_37_active;
  logic stage_38_active;
  logic stage_39_active;
  logic stage_40_active;
  logic stage_41_active;
  logic stage_42_active;
  logic stage_43_active;
  logic stage_44_active;
  logic stage_45_active;
  logic stage_46_active;
  logic stage_47_active;
  logic stage_48_active;
  logic stage_49_active;
  logic stage_50_active;
  logic stage_51_active;
  logic stage_52_active;
  logic stage_53_active;
  logic stage_54_active;
  logic stage_55_active;
  logic stage_56_active;
  logic stage_57_active;
  logic stage_58_active;
  logic stage_59_active;
  logic stage_60_active;
  logic stage_61_active;
  logic stage_62_active;
  logic stage_63_active;
  logic stage_64_active;
  logic stage_65_active;
  logic stage_66_active;
  logic stage_67_active;
  logic stage_68_active;
  logic stage_69_active;
  logic stage_70_active;
  logic stage_71_active;
  logic stage_72_active;
  logic stage_73_active;
  logic stage_74_active;
  logic stage_75_active;
  logic stage_76_active;
  logic stage_77_active;
  logic stage_78_active;
  logic stage_79_active;
  logic stage_80_active;
  logic stage_81_active;
  logic stage_82_active;
  logic stage_83_active;
  logic stage_84_active;
  logic stage_85_active;
  logic stage_86_active;
  logic stage_87_active;
  logic stage_88_active;
  logic stage_89_active;
  logic stage_90_active;
  logic stage_91_active;
  logic stage_92_active;
  logic stage_93_active;
  logic stage_94_active;
  logic stage_95_active;
  logic stage_96_active;
  logic stage_97_active;
  logic stage_98_active;
  logic stage_99_active;
  logic stage_100_active;
  logic stage_101_active;
  logic stage_102_active;
  logic stage_103_active;
  logic stage_104_active;
  logic stage_105_active;
  logic stage_106_active;
  logic stage_107_active;
  logic stage_108_active;
  logic stage_109_active;
  logic stage_110_active;
  logic stage_111_active;
  logic stage_112_active;
  logic stage_113_active;
  logic stage_114_active;
  logic stage_115_active;
  logic stage_116_active;
  logic stage_117_active;
  logic stage_118_active;
  logic stage_119_active;
  logic stage_120_active;
  logic stage_121_active;
  logic stage_122_active;
  logic stage_123_active;
  logic stage_124_active;
  logic stage_125_active;
  logic stage_126_active;
  logic stage_127_active;
  logic stage_128_active;
  logic stage_129_active;
  logic stage_130_active;
  logic stage_131_active;
  logic stage_132_active;
  logic stage_133_active;
  logic stage_134_active;
  logic stage_135_active;
  logic stage_136_active;
  logic stage_137_active;
  logic stage_138_active;
  logic stage_139_active;
  logic stage_140_active;
  logic stage_141_active;
  logic stage_142_active;
  logic stage_143_active;
  logic stage_144_active;
  logic stage_145_active;
  logic stage_146_active;
  logic stage_147_active;
  logic stage_148_active;
  logic stage_149_active;
  logic stage_150_active;
  logic stage_151_active;
  logic stage_152_active;
  logic stage_153_active;
  logic stage_154_active;
  logic stage_155_active;
  logic stage_156_active;
  logic stage_157_active;
  logic stage_158_active;
  logic stage_159_active;
  logic stage_160_active;
  logic stage_161_active;
  logic stage_162_active;
  logic stage_163_active;
  logic stage_164_active;
  logic stage_165_active;
  logic stage_166_active;
  logic stage_167_active;
  logic stage_168_active;
  logic stage_169_active;
  logic stage_170_active;
  logic stage_171_active;
  logic stage_172_active;
  logic stage_173_active;
  logic stage_174_active;
  logic stage_175_active;
  logic stage_176_active;
  logic stage_177_active;
  logic stage_178_active;
  logic stage_179_active;
  logic stage_180_active;

  logic stage_0_at_iter_0;
  logic stage_1_at_iter_0;
  logic stage_2_at_iter_0;
  logic stage_3_at_iter_0;
  logic stage_4_at_iter_0;
  logic stage_5_at_iter_0;
  logic stage_6_at_iter_0;
  logic stage_7_at_iter_0;
  logic stage_8_at_iter_0;
  logic stage_9_at_iter_0;
  logic stage_10_at_iter_0;
  logic stage_11_at_iter_0;
  logic stage_12_at_iter_0;
  logic stage_13_at_iter_0;
  logic stage_14_at_iter_0;
  logic stage_15_at_iter_0;
  logic stage_16_at_iter_0;
  logic stage_17_at_iter_0;
  logic stage_18_at_iter_0;
  logic stage_19_at_iter_0;
  logic stage_20_at_iter_0;
  logic stage_21_at_iter_0;
  logic stage_22_at_iter_0;
  logic stage_23_at_iter_0;
  logic stage_24_at_iter_0;
  logic stage_25_at_iter_0;
  logic stage_26_at_iter_0;
  logic stage_27_at_iter_0;
  logic stage_28_at_iter_0;
  logic stage_29_at_iter_0;
  logic stage_30_at_iter_0;
  logic stage_31_at_iter_0;
  logic stage_32_at_iter_0;
  logic stage_33_at_iter_0;
  logic stage_34_at_iter_0;
  logic stage_35_at_iter_0;
  logic stage_36_at_iter_0;
  logic stage_37_at_iter_0;
  logic stage_38_at_iter_0;
  logic stage_39_at_iter_0;
  logic stage_40_at_iter_0;
  logic stage_41_at_iter_0;
  logic stage_42_at_iter_0;
  logic stage_43_at_iter_0;
  logic stage_44_at_iter_0;
  logic stage_45_at_iter_0;
  logic stage_46_at_iter_0;
  logic stage_47_at_iter_0;
  logic stage_48_at_iter_0;
  logic stage_49_at_iter_0;
  logic stage_50_at_iter_0;
  logic stage_51_at_iter_0;
  logic stage_52_at_iter_0;
  logic stage_53_at_iter_0;
  logic stage_54_at_iter_0;
  logic stage_55_at_iter_0;
  logic stage_56_at_iter_0;
  logic stage_57_at_iter_0;
  logic stage_58_at_iter_0;
  logic stage_59_at_iter_0;
  logic stage_60_at_iter_0;
  logic stage_61_at_iter_0;
  logic stage_62_at_iter_0;
  logic stage_63_at_iter_0;
  logic stage_64_at_iter_0;
  logic stage_65_at_iter_0;
  logic stage_66_at_iter_0;
  logic stage_67_at_iter_0;
  logic stage_68_at_iter_0;
  logic stage_69_at_iter_0;
  logic stage_70_at_iter_0;
  logic stage_71_at_iter_0;
  logic stage_72_at_iter_0;
  logic stage_73_at_iter_0;
  logic stage_74_at_iter_0;
  logic stage_75_at_iter_0;
  logic stage_76_at_iter_0;
  logic stage_77_at_iter_0;
  logic stage_78_at_iter_0;
  logic stage_79_at_iter_0;
  logic stage_80_at_iter_0;
  logic stage_81_at_iter_0;
  logic stage_82_at_iter_0;
  logic stage_83_at_iter_0;
  logic stage_84_at_iter_0;
  logic stage_85_at_iter_0;
  logic stage_86_at_iter_0;
  logic stage_87_at_iter_0;
  logic stage_88_at_iter_0;
  logic stage_89_at_iter_0;
  logic stage_90_at_iter_0;
  logic stage_91_at_iter_0;
  logic stage_92_at_iter_0;
  logic stage_93_at_iter_0;
  logic stage_94_at_iter_0;
  logic stage_95_at_iter_0;
  logic stage_96_at_iter_0;
  logic stage_97_at_iter_0;
  logic stage_98_at_iter_0;
  logic stage_99_at_iter_0;
  logic stage_100_at_iter_0;
  logic stage_101_at_iter_0;
  logic stage_102_at_iter_0;
  logic stage_103_at_iter_0;
  logic stage_104_at_iter_0;
  logic stage_105_at_iter_0;
  logic stage_106_at_iter_0;
  logic stage_107_at_iter_0;
  logic stage_108_at_iter_0;
  logic stage_109_at_iter_0;
  logic stage_110_at_iter_0;
  logic stage_111_at_iter_0;
  logic stage_112_at_iter_0;
  logic stage_113_at_iter_0;
  logic stage_114_at_iter_0;
  logic stage_115_at_iter_0;
  logic stage_116_at_iter_0;
  logic stage_117_at_iter_0;
  logic stage_118_at_iter_0;
  logic stage_119_at_iter_0;
  logic stage_120_at_iter_0;
  logic stage_121_at_iter_0;
  logic stage_122_at_iter_0;
  logic stage_123_at_iter_0;
  logic stage_124_at_iter_0;
  logic stage_125_at_iter_0;
  logic stage_126_at_iter_0;
  logic stage_127_at_iter_0;
  logic stage_128_at_iter_0;
  logic stage_129_at_iter_0;
  logic stage_130_at_iter_0;
  logic stage_131_at_iter_0;
  logic stage_132_at_iter_0;
  logic stage_133_at_iter_0;
  logic stage_134_at_iter_0;
  logic stage_135_at_iter_0;
  logic stage_136_at_iter_0;
  logic stage_137_at_iter_0;
  logic stage_138_at_iter_0;
  logic stage_139_at_iter_0;
  logic stage_140_at_iter_0;
  logic stage_141_at_iter_0;
  logic stage_142_at_iter_0;
  logic stage_143_at_iter_0;
  logic stage_144_at_iter_0;
  logic stage_145_at_iter_0;
  logic stage_146_at_iter_0;
  logic stage_147_at_iter_0;
  logic stage_148_at_iter_0;
  logic stage_149_at_iter_0;
  logic stage_150_at_iter_0;
  logic stage_151_at_iter_0;
  logic stage_152_at_iter_0;
  logic stage_153_at_iter_0;
  logic stage_154_at_iter_0;
  logic stage_155_at_iter_0;
  logic stage_156_at_iter_0;
  logic stage_157_at_iter_0;
  logic stage_158_at_iter_0;
  logic stage_159_at_iter_0;
  logic stage_160_at_iter_0;
  logic stage_161_at_iter_0;
  logic stage_162_at_iter_0;
  logic stage_163_at_iter_0;
  logic stage_164_at_iter_0;
  logic stage_165_at_iter_0;
  logic stage_166_at_iter_0;
  logic stage_167_at_iter_0;
  logic stage_168_at_iter_0;
  logic stage_169_at_iter_0;
  logic stage_170_at_iter_0;
  logic stage_171_at_iter_0;
  logic stage_172_at_iter_0;
  logic stage_173_at_iter_0;
  logic stage_174_at_iter_0;
  logic stage_175_at_iter_0;
  logic stage_176_at_iter_0;
  logic stage_177_at_iter_0;
  logic stage_178_at_iter_0;
  logic stage_179_at_iter_0;
  logic stage_180_at_iter_0;

  assign stage_0_active = start | started;
  assign stage_0_at_iter_0 = start;
  assign done = stage_180_active;

  // Pipeline datapath registers...
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_2;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_3;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_4;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_5;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_6;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_7;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_8;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_9;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_10;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_11;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_12;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_13;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_14;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_15;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_16;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_17;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_18;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_19;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_20;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_21;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_22;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_23;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_24;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_25;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_26;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_27;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_28;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_29;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_30;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_31;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_32;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_33;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_34;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_35;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_36;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_37;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_38;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_39;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_40;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_41;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_42;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_43;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_44;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_45;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_46;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_47;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_48;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_49;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_50;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_51;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_52;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_53;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_54;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_55;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_56;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_57;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_58;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_59;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_60;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_61;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_62;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_63;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_64;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_65;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_66;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_67;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_68;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_69;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_70;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_71;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_72;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_73;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_74;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_75;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_76;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_77;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_78;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_79;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_80;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_81;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_82;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_83;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_84;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_85;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_86;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_87;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_88;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_89;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_90;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_91;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_92;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_93;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_94;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_95;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_96;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_97;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_98;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_99;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_100;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_101;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_102;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_103;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_104;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_105;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_106;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_107;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_108;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_109;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_110;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_111;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_112;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_113;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_114;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_115;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_116;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_117;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_118;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_119;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_120;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_121;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_122;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_123;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_124;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_125;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_126;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_127;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_128;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_129;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_130;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_131;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_132;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_133;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_134;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_135;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_136;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_137;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_138;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_139;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_140;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_141;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_142;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_143;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_144;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_145;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_146;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_147;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_148;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_149;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_150;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_151;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_152;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_153;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_154;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_155;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_156;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_157;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_158;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_159;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_160;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_161;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_162;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_163;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_164;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_165;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_166;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_167;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_168;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_169;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_170;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_171;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_172;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_173;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_174;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_175;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_176;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_177;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_178;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_179;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_180;
  reg [31:0] in_off_chip_in_update_0_read_read_0_stage_181;
  reg [31:0] in_update_0_stage_3;
  reg [31:0] in_update_0_stage_4;
  reg [31:0] in_update_0_stage_5;
  reg [31:0] in_update_0_stage_6;
  reg [31:0] in_update_0_stage_7;
  reg [31:0] in_update_0_stage_8;
  reg [31:0] in_update_0_stage_9;
  reg [31:0] in_update_0_stage_10;
  reg [31:0] in_update_0_stage_11;
  reg [31:0] in_update_0_stage_12;
  reg [31:0] in_update_0_stage_13;
  reg [31:0] in_update_0_stage_14;
  reg [31:0] in_update_0_stage_15;
  reg [31:0] in_update_0_stage_16;
  reg [31:0] in_update_0_stage_17;
  reg [31:0] in_update_0_stage_18;
  reg [31:0] in_update_0_stage_19;
  reg [31:0] in_update_0_stage_20;
  reg [31:0] in_update_0_stage_21;
  reg [31:0] in_update_0_stage_22;
  reg [31:0] in_update_0_stage_23;
  reg [31:0] in_update_0_stage_24;
  reg [31:0] in_update_0_stage_25;
  reg [31:0] in_update_0_stage_26;
  reg [31:0] in_update_0_stage_27;
  reg [31:0] in_update_0_stage_28;
  reg [31:0] in_update_0_stage_29;
  reg [31:0] in_update_0_stage_30;
  reg [31:0] in_update_0_stage_31;
  reg [31:0] in_update_0_stage_32;
  reg [31:0] in_update_0_stage_33;
  reg [31:0] in_update_0_stage_34;
  reg [31:0] in_update_0_stage_35;
  reg [31:0] in_update_0_stage_36;
  reg [31:0] in_update_0_stage_37;
  reg [31:0] in_update_0_stage_38;
  reg [31:0] in_update_0_stage_39;
  reg [31:0] in_update_0_stage_40;
  reg [31:0] in_update_0_stage_41;
  reg [31:0] in_update_0_stage_42;
  reg [31:0] in_update_0_stage_43;
  reg [31:0] in_update_0_stage_44;
  reg [31:0] in_update_0_stage_45;
  reg [31:0] in_update_0_stage_46;
  reg [31:0] in_update_0_stage_47;
  reg [31:0] in_update_0_stage_48;
  reg [31:0] in_update_0_stage_49;
  reg [31:0] in_update_0_stage_50;
  reg [31:0] in_update_0_stage_51;
  reg [31:0] in_update_0_stage_52;
  reg [31:0] in_update_0_stage_53;
  reg [31:0] in_update_0_stage_54;
  reg [31:0] in_update_0_stage_55;
  reg [31:0] in_update_0_stage_56;
  reg [31:0] in_update_0_stage_57;
  reg [31:0] in_update_0_stage_58;
  reg [31:0] in_update_0_stage_59;
  reg [31:0] in_update_0_stage_60;
  reg [31:0] in_update_0_stage_61;
  reg [31:0] in_update_0_stage_62;
  reg [31:0] in_update_0_stage_63;
  reg [31:0] in_update_0_stage_64;
  reg [31:0] in_update_0_stage_65;
  reg [31:0] in_update_0_stage_66;
  reg [31:0] in_update_0_stage_67;
  reg [31:0] in_update_0_stage_68;
  reg [31:0] in_update_0_stage_69;
  reg [31:0] in_update_0_stage_70;
  reg [31:0] in_update_0_stage_71;
  reg [31:0] in_update_0_stage_72;
  reg [31:0] in_update_0_stage_73;
  reg [31:0] in_update_0_stage_74;
  reg [31:0] in_update_0_stage_75;
  reg [31:0] in_update_0_stage_76;
  reg [31:0] in_update_0_stage_77;
  reg [31:0] in_update_0_stage_78;
  reg [31:0] in_update_0_stage_79;
  reg [31:0] in_update_0_stage_80;
  reg [31:0] in_update_0_stage_81;
  reg [31:0] in_update_0_stage_82;
  reg [31:0] in_update_0_stage_83;
  reg [31:0] in_update_0_stage_84;
  reg [31:0] in_update_0_stage_85;
  reg [31:0] in_update_0_stage_86;
  reg [31:0] in_update_0_stage_87;
  reg [31:0] in_update_0_stage_88;
  reg [31:0] in_update_0_stage_89;
  reg [31:0] in_update_0_stage_90;
  reg [31:0] in_update_0_stage_91;
  reg [31:0] in_update_0_stage_92;
  reg [31:0] in_update_0_stage_93;
  reg [31:0] in_update_0_stage_94;
  reg [31:0] in_update_0_stage_95;
  reg [31:0] in_update_0_stage_96;
  reg [31:0] in_update_0_stage_97;
  reg [31:0] in_update_0_stage_98;
  reg [31:0] in_update_0_stage_99;
  reg [31:0] in_update_0_stage_100;
  reg [31:0] in_update_0_stage_101;
  reg [31:0] in_update_0_stage_102;
  reg [31:0] in_update_0_stage_103;
  reg [31:0] in_update_0_stage_104;
  reg [31:0] in_update_0_stage_105;
  reg [31:0] in_update_0_stage_106;
  reg [31:0] in_update_0_stage_107;
  reg [31:0] in_update_0_stage_108;
  reg [31:0] in_update_0_stage_109;
  reg [31:0] in_update_0_stage_110;
  reg [31:0] in_update_0_stage_111;
  reg [31:0] in_update_0_stage_112;
  reg [31:0] in_update_0_stage_113;
  reg [31:0] in_update_0_stage_114;
  reg [31:0] in_update_0_stage_115;
  reg [31:0] in_update_0_stage_116;
  reg [31:0] in_update_0_stage_117;
  reg [31:0] in_update_0_stage_118;
  reg [31:0] in_update_0_stage_119;
  reg [31:0] in_update_0_stage_120;
  reg [31:0] in_update_0_stage_121;
  reg [31:0] in_update_0_stage_122;
  reg [31:0] in_update_0_stage_123;
  reg [31:0] in_update_0_stage_124;
  reg [31:0] in_update_0_stage_125;
  reg [31:0] in_update_0_stage_126;
  reg [31:0] in_update_0_stage_127;
  reg [31:0] in_update_0_stage_128;
  reg [31:0] in_update_0_stage_129;
  reg [31:0] in_update_0_stage_130;
  reg [31:0] in_update_0_stage_131;
  reg [31:0] in_update_0_stage_132;
  reg [31:0] in_update_0_stage_133;
  reg [31:0] in_update_0_stage_134;
  reg [31:0] in_update_0_stage_135;
  reg [31:0] in_update_0_stage_136;
  reg [31:0] in_update_0_stage_137;
  reg [31:0] in_update_0_stage_138;
  reg [31:0] in_update_0_stage_139;
  reg [31:0] in_update_0_stage_140;
  reg [31:0] in_update_0_stage_141;
  reg [31:0] in_update_0_stage_142;
  reg [31:0] in_update_0_stage_143;
  reg [31:0] in_update_0_stage_144;
  reg [31:0] in_update_0_stage_145;
  reg [31:0] in_update_0_stage_146;
  reg [31:0] in_update_0_stage_147;
  reg [31:0] in_update_0_stage_148;
  reg [31:0] in_update_0_stage_149;
  reg [31:0] in_update_0_stage_150;
  reg [31:0] in_update_0_stage_151;
  reg [31:0] in_update_0_stage_152;
  reg [31:0] in_update_0_stage_153;
  reg [31:0] in_update_0_stage_154;
  reg [31:0] in_update_0_stage_155;
  reg [31:0] in_update_0_stage_156;
  reg [31:0] in_update_0_stage_157;
  reg [31:0] in_update_0_stage_158;
  reg [31:0] in_update_0_stage_159;
  reg [31:0] in_update_0_stage_160;
  reg [31:0] in_update_0_stage_161;
  reg [31:0] in_update_0_stage_162;
  reg [31:0] in_update_0_stage_163;
  reg [31:0] in_update_0_stage_164;
  reg [31:0] in_update_0_stage_165;
  reg [31:0] in_update_0_stage_166;
  reg [31:0] in_update_0_stage_167;
  reg [31:0] in_update_0_stage_168;
  reg [31:0] in_update_0_stage_169;
  reg [31:0] in_update_0_stage_170;
  reg [31:0] in_update_0_stage_171;
  reg [31:0] in_update_0_stage_172;
  reg [31:0] in_update_0_stage_173;
  reg [31:0] in_update_0_stage_174;
  reg [31:0] in_update_0_stage_175;
  reg [31:0] in_update_0_stage_176;
  reg [31:0] in_update_0_stage_177;
  reg [31:0] in_update_0_stage_178;
  reg [31:0] in_update_0_stage_179;
  reg [31:0] in_update_0_stage_180;
  reg [31:0] in_update_0_stage_181;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_8;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_9;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_10;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_11;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_12;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_13;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_14;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_15;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_16;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_17;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_18;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_19;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_20;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_21;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_22;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_23;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_24;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_25;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_26;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_27;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_28;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_29;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_30;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_31;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_32;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_33;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_34;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_35;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_36;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_37;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_38;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_39;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_40;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_41;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_42;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_43;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_44;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_45;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_46;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_47;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_48;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_49;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_50;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_51;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_52;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_53;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_54;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_55;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_56;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_57;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_58;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_59;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_60;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_61;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_62;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_63;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_64;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_65;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_66;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_67;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_68;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_69;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_70;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_71;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_72;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_73;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_74;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_75;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_76;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_77;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_78;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_79;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_80;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_81;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_82;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_83;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_84;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_85;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_86;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_87;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_88;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_89;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_90;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_91;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_92;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_93;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_94;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_95;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_96;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_97;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_98;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_99;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_100;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_101;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_102;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_103;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_104;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_105;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_106;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_107;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_108;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_109;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_110;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_111;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_112;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_113;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_114;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_115;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_116;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_117;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_118;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_119;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_120;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_121;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_122;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_123;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_124;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_125;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_126;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_127;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_128;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_129;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_130;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_131;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_132;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_133;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_134;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_135;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_136;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_137;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_138;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_139;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_140;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_141;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_142;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_143;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_144;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_145;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_146;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_147;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_148;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_149;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_150;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_151;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_152;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_153;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_154;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_155;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_156;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_157;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_158;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_159;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_160;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_161;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_162;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_163;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_164;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_165;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_166;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_167;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_168;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_169;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_170;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_171;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_172;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_173;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_174;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_175;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_176;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_177;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_178;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_179;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_180;
  reg [31:0] bright_bright_weights_update_0_read_read_4_stage_181;
  reg [31:0] bright_weights_update_0_stage_9;
  reg [31:0] bright_weights_update_0_stage_10;
  reg [31:0] bright_weights_update_0_stage_11;
  reg [31:0] bright_weights_update_0_stage_12;
  reg [31:0] bright_weights_update_0_stage_13;
  reg [31:0] bright_weights_update_0_stage_14;
  reg [31:0] bright_weights_update_0_stage_15;
  reg [31:0] bright_weights_update_0_stage_16;
  reg [31:0] bright_weights_update_0_stage_17;
  reg [31:0] bright_weights_update_0_stage_18;
  reg [31:0] bright_weights_update_0_stage_19;
  reg [31:0] bright_weights_update_0_stage_20;
  reg [31:0] bright_weights_update_0_stage_21;
  reg [31:0] bright_weights_update_0_stage_22;
  reg [31:0] bright_weights_update_0_stage_23;
  reg [31:0] bright_weights_update_0_stage_24;
  reg [31:0] bright_weights_update_0_stage_25;
  reg [31:0] bright_weights_update_0_stage_26;
  reg [31:0] bright_weights_update_0_stage_27;
  reg [31:0] bright_weights_update_0_stage_28;
  reg [31:0] bright_weights_update_0_stage_29;
  reg [31:0] bright_weights_update_0_stage_30;
  reg [31:0] bright_weights_update_0_stage_31;
  reg [31:0] bright_weights_update_0_stage_32;
  reg [31:0] bright_weights_update_0_stage_33;
  reg [31:0] bright_weights_update_0_stage_34;
  reg [31:0] bright_weights_update_0_stage_35;
  reg [31:0] bright_weights_update_0_stage_36;
  reg [31:0] bright_weights_update_0_stage_37;
  reg [31:0] bright_weights_update_0_stage_38;
  reg [31:0] bright_weights_update_0_stage_39;
  reg [31:0] bright_weights_update_0_stage_40;
  reg [31:0] bright_weights_update_0_stage_41;
  reg [31:0] bright_weights_update_0_stage_42;
  reg [31:0] bright_weights_update_0_stage_43;
  reg [31:0] bright_weights_update_0_stage_44;
  reg [31:0] bright_weights_update_0_stage_45;
  reg [31:0] bright_weights_update_0_stage_46;
  reg [31:0] bright_weights_update_0_stage_47;
  reg [31:0] bright_weights_update_0_stage_48;
  reg [31:0] bright_weights_update_0_stage_49;
  reg [31:0] bright_weights_update_0_stage_50;
  reg [31:0] bright_weights_update_0_stage_51;
  reg [31:0] bright_weights_update_0_stage_52;
  reg [31:0] bright_weights_update_0_stage_53;
  reg [31:0] bright_weights_update_0_stage_54;
  reg [31:0] bright_weights_update_0_stage_55;
  reg [31:0] bright_weights_update_0_stage_56;
  reg [31:0] bright_weights_update_0_stage_57;
  reg [31:0] bright_weights_update_0_stage_58;
  reg [31:0] bright_weights_update_0_stage_59;
  reg [31:0] bright_weights_update_0_stage_60;
  reg [31:0] bright_weights_update_0_stage_61;
  reg [31:0] bright_weights_update_0_stage_62;
  reg [31:0] bright_weights_update_0_stage_63;
  reg [31:0] bright_weights_update_0_stage_64;
  reg [31:0] bright_weights_update_0_stage_65;
  reg [31:0] bright_weights_update_0_stage_66;
  reg [31:0] bright_weights_update_0_stage_67;
  reg [31:0] bright_weights_update_0_stage_68;
  reg [31:0] bright_weights_update_0_stage_69;
  reg [31:0] bright_weights_update_0_stage_70;
  reg [31:0] bright_weights_update_0_stage_71;
  reg [31:0] bright_weights_update_0_stage_72;
  reg [31:0] bright_weights_update_0_stage_73;
  reg [31:0] bright_weights_update_0_stage_74;
  reg [31:0] bright_weights_update_0_stage_75;
  reg [31:0] bright_weights_update_0_stage_76;
  reg [31:0] bright_weights_update_0_stage_77;
  reg [31:0] bright_weights_update_0_stage_78;
  reg [31:0] bright_weights_update_0_stage_79;
  reg [31:0] bright_weights_update_0_stage_80;
  reg [31:0] bright_weights_update_0_stage_81;
  reg [31:0] bright_weights_update_0_stage_82;
  reg [31:0] bright_weights_update_0_stage_83;
  reg [31:0] bright_weights_update_0_stage_84;
  reg [31:0] bright_weights_update_0_stage_85;
  reg [31:0] bright_weights_update_0_stage_86;
  reg [31:0] bright_weights_update_0_stage_87;
  reg [31:0] bright_weights_update_0_stage_88;
  reg [31:0] bright_weights_update_0_stage_89;
  reg [31:0] bright_weights_update_0_stage_90;
  reg [31:0] bright_weights_update_0_stage_91;
  reg [31:0] bright_weights_update_0_stage_92;
  reg [31:0] bright_weights_update_0_stage_93;
  reg [31:0] bright_weights_update_0_stage_94;
  reg [31:0] bright_weights_update_0_stage_95;
  reg [31:0] bright_weights_update_0_stage_96;
  reg [31:0] bright_weights_update_0_stage_97;
  reg [31:0] bright_weights_update_0_stage_98;
  reg [31:0] bright_weights_update_0_stage_99;
  reg [31:0] bright_weights_update_0_stage_100;
  reg [31:0] bright_weights_update_0_stage_101;
  reg [31:0] bright_weights_update_0_stage_102;
  reg [31:0] bright_weights_update_0_stage_103;
  reg [31:0] bright_weights_update_0_stage_104;
  reg [31:0] bright_weights_update_0_stage_105;
  reg [31:0] bright_weights_update_0_stage_106;
  reg [31:0] bright_weights_update_0_stage_107;
  reg [31:0] bright_weights_update_0_stage_108;
  reg [31:0] bright_weights_update_0_stage_109;
  reg [31:0] bright_weights_update_0_stage_110;
  reg [31:0] bright_weights_update_0_stage_111;
  reg [31:0] bright_weights_update_0_stage_112;
  reg [31:0] bright_weights_update_0_stage_113;
  reg [31:0] bright_weights_update_0_stage_114;
  reg [31:0] bright_weights_update_0_stage_115;
  reg [31:0] bright_weights_update_0_stage_116;
  reg [31:0] bright_weights_update_0_stage_117;
  reg [31:0] bright_weights_update_0_stage_118;
  reg [31:0] bright_weights_update_0_stage_119;
  reg [31:0] bright_weights_update_0_stage_120;
  reg [31:0] bright_weights_update_0_stage_121;
  reg [31:0] bright_weights_update_0_stage_122;
  reg [31:0] bright_weights_update_0_stage_123;
  reg [31:0] bright_weights_update_0_stage_124;
  reg [31:0] bright_weights_update_0_stage_125;
  reg [31:0] bright_weights_update_0_stage_126;
  reg [31:0] bright_weights_update_0_stage_127;
  reg [31:0] bright_weights_update_0_stage_128;
  reg [31:0] bright_weights_update_0_stage_129;
  reg [31:0] bright_weights_update_0_stage_130;
  reg [31:0] bright_weights_update_0_stage_131;
  reg [31:0] bright_weights_update_0_stage_132;
  reg [31:0] bright_weights_update_0_stage_133;
  reg [31:0] bright_weights_update_0_stage_134;
  reg [31:0] bright_weights_update_0_stage_135;
  reg [31:0] bright_weights_update_0_stage_136;
  reg [31:0] bright_weights_update_0_stage_137;
  reg [31:0] bright_weights_update_0_stage_138;
  reg [31:0] bright_weights_update_0_stage_139;
  reg [31:0] bright_weights_update_0_stage_140;
  reg [31:0] bright_weights_update_0_stage_141;
  reg [31:0] bright_weights_update_0_stage_142;
  reg [31:0] bright_weights_update_0_stage_143;
  reg [31:0] bright_weights_update_0_stage_144;
  reg [31:0] bright_weights_update_0_stage_145;
  reg [31:0] bright_weights_update_0_stage_146;
  reg [31:0] bright_weights_update_0_stage_147;
  reg [31:0] bright_weights_update_0_stage_148;
  reg [31:0] bright_weights_update_0_stage_149;
  reg [31:0] bright_weights_update_0_stage_150;
  reg [31:0] bright_weights_update_0_stage_151;
  reg [31:0] bright_weights_update_0_stage_152;
  reg [31:0] bright_weights_update_0_stage_153;
  reg [31:0] bright_weights_update_0_stage_154;
  reg [31:0] bright_weights_update_0_stage_155;
  reg [31:0] bright_weights_update_0_stage_156;
  reg [31:0] bright_weights_update_0_stage_157;
  reg [31:0] bright_weights_update_0_stage_158;
  reg [31:0] bright_weights_update_0_stage_159;
  reg [31:0] bright_weights_update_0_stage_160;
  reg [31:0] bright_weights_update_0_stage_161;
  reg [31:0] bright_weights_update_0_stage_162;
  reg [31:0] bright_weights_update_0_stage_163;
  reg [31:0] bright_weights_update_0_stage_164;
  reg [31:0] bright_weights_update_0_stage_165;
  reg [31:0] bright_weights_update_0_stage_166;
  reg [31:0] bright_weights_update_0_stage_167;
  reg [31:0] bright_weights_update_0_stage_168;
  reg [31:0] bright_weights_update_0_stage_169;
  reg [31:0] bright_weights_update_0_stage_170;
  reg [31:0] bright_weights_update_0_stage_171;
  reg [31:0] bright_weights_update_0_stage_172;
  reg [31:0] bright_weights_update_0_stage_173;
  reg [31:0] bright_weights_update_0_stage_174;
  reg [31:0] bright_weights_update_0_stage_175;
  reg [31:0] bright_weights_update_0_stage_176;
  reg [31:0] bright_weights_update_0_stage_177;
  reg [31:0] bright_weights_update_0_stage_178;
  reg [31:0] bright_weights_update_0_stage_179;
  reg [31:0] bright_weights_update_0_stage_180;
  reg [31:0] bright_weights_update_0_stage_181;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_10;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_11;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_12;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_13;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_14;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_15;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_16;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_17;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_18;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_19;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_20;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_21;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_22;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_23;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_24;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_25;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_26;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_27;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_28;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_29;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_30;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_31;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_32;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_33;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_34;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_35;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_36;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_37;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_38;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_39;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_40;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_41;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_42;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_43;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_44;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_45;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_46;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_47;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_48;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_49;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_50;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_51;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_52;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_53;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_54;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_55;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_56;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_57;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_58;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_59;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_60;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_61;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_62;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_63;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_64;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_65;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_66;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_67;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_68;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_69;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_70;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_71;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_72;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_73;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_74;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_75;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_76;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_77;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_78;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_79;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_80;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_81;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_82;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_83;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_84;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_85;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_86;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_87;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_88;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_89;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_90;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_91;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_92;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_93;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_94;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_95;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_96;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_97;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_98;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_99;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_100;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_101;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_102;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_103;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_104;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_105;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_106;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_107;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_108;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_109;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_110;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_111;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_112;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_113;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_114;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_115;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_116;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_117;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_118;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_119;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_120;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_121;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_122;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_123;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_124;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_125;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_126;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_127;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_128;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_129;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_130;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_131;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_132;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_133;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_134;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_135;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_136;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_137;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_138;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_139;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_140;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_141;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_142;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_143;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_144;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_145;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_146;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_147;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_148;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_149;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_150;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_151;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_152;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_153;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_154;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_155;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_156;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_157;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_158;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_159;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_160;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_161;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_162;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_163;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_164;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_165;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_166;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_167;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_168;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_169;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_170;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_171;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_172;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_173;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_174;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_175;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_176;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_177;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_178;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_179;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_180;
  reg [31:0] bright_weights_bright_weights_update_0_write_write_5_stage_181;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_85;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_86;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_87;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_88;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_89;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_90;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_91;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_92;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_93;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_94;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_95;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_96;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_97;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_98;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_99;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_100;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_101;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_102;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_103;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_104;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_105;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_106;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_107;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_108;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_109;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_110;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_111;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_112;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_113;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_114;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_115;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_116;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_117;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_118;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_119;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_120;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_121;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_122;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_123;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_124;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_125;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_126;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_127;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_128;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_129;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_130;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_131;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_132;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_133;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_134;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_135;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_136;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_137;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_138;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_139;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_140;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_141;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_142;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_143;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_144;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_145;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_146;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_147;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_148;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_149;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_150;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_151;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_152;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_153;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_154;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_155;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_156;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_157;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_158;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_159;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_160;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_161;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_162;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_163;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_164;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_165;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_166;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_167;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_168;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_169;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_170;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_171;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_172;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_173;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_174;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_175;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_176;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_177;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_178;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_179;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_180;
  reg [287:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_181;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_14;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_15;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_16;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_17;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_18;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_19;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_20;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_21;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_22;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_23;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_24;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_25;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_26;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_27;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_28;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_29;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_30;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_31;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_32;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_33;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_34;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_35;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_36;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_37;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_38;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_39;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_40;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_41;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_42;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_43;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_44;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_45;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_46;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_47;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_48;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_49;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_50;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_51;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_52;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_53;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_54;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_55;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_56;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_57;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_58;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_59;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_60;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_61;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_62;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_63;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_64;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_65;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_66;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_67;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_68;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_69;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_70;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_71;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_72;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_73;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_74;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_75;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_76;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_77;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_78;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_79;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_80;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_81;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_82;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_83;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_84;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_85;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_86;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_87;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_88;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_89;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_90;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_91;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_92;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_93;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_94;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_95;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_96;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_97;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_98;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_99;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_100;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_101;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_102;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_103;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_104;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_105;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_106;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_107;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_108;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_109;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_110;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_111;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_112;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_113;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_114;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_115;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_116;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_117;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_118;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_119;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_120;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_121;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_122;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_123;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_124;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_125;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_126;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_127;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_128;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_129;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_130;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_131;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_132;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_133;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_134;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_135;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_136;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_137;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_138;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_139;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_140;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_141;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_142;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_143;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_144;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_145;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_146;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_147;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_148;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_149;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_150;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_151;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_152;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_153;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_154;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_155;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_156;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_157;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_158;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_159;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_160;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_161;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_162;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_163;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_164;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_165;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_166;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_167;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_168;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_169;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_170;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_171;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_172;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_173;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_174;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_175;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_176;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_177;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_178;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_179;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_180;
  reg [31:0] dark_dark_weights_update_0_read_read_8_stage_181;
  reg [31:0] dark_weights_update_0_stage_15;
  reg [31:0] dark_weights_update_0_stage_16;
  reg [31:0] dark_weights_update_0_stage_17;
  reg [31:0] dark_weights_update_0_stage_18;
  reg [31:0] dark_weights_update_0_stage_19;
  reg [31:0] dark_weights_update_0_stage_20;
  reg [31:0] dark_weights_update_0_stage_21;
  reg [31:0] dark_weights_update_0_stage_22;
  reg [31:0] dark_weights_update_0_stage_23;
  reg [31:0] dark_weights_update_0_stage_24;
  reg [31:0] dark_weights_update_0_stage_25;
  reg [31:0] dark_weights_update_0_stage_26;
  reg [31:0] dark_weights_update_0_stage_27;
  reg [31:0] dark_weights_update_0_stage_28;
  reg [31:0] dark_weights_update_0_stage_29;
  reg [31:0] dark_weights_update_0_stage_30;
  reg [31:0] dark_weights_update_0_stage_31;
  reg [31:0] dark_weights_update_0_stage_32;
  reg [31:0] dark_weights_update_0_stage_33;
  reg [31:0] dark_weights_update_0_stage_34;
  reg [31:0] dark_weights_update_0_stage_35;
  reg [31:0] dark_weights_update_0_stage_36;
  reg [31:0] dark_weights_update_0_stage_37;
  reg [31:0] dark_weights_update_0_stage_38;
  reg [31:0] dark_weights_update_0_stage_39;
  reg [31:0] dark_weights_update_0_stage_40;
  reg [31:0] dark_weights_update_0_stage_41;
  reg [31:0] dark_weights_update_0_stage_42;
  reg [31:0] dark_weights_update_0_stage_43;
  reg [31:0] dark_weights_update_0_stage_44;
  reg [31:0] dark_weights_update_0_stage_45;
  reg [31:0] dark_weights_update_0_stage_46;
  reg [31:0] dark_weights_update_0_stage_47;
  reg [31:0] dark_weights_update_0_stage_48;
  reg [31:0] dark_weights_update_0_stage_49;
  reg [31:0] dark_weights_update_0_stage_50;
  reg [31:0] dark_weights_update_0_stage_51;
  reg [31:0] dark_weights_update_0_stage_52;
  reg [31:0] dark_weights_update_0_stage_53;
  reg [31:0] dark_weights_update_0_stage_54;
  reg [31:0] dark_weights_update_0_stage_55;
  reg [31:0] dark_weights_update_0_stage_56;
  reg [31:0] dark_weights_update_0_stage_57;
  reg [31:0] dark_weights_update_0_stage_58;
  reg [31:0] dark_weights_update_0_stage_59;
  reg [31:0] dark_weights_update_0_stage_60;
  reg [31:0] dark_weights_update_0_stage_61;
  reg [31:0] dark_weights_update_0_stage_62;
  reg [31:0] dark_weights_update_0_stage_63;
  reg [31:0] dark_weights_update_0_stage_64;
  reg [31:0] dark_weights_update_0_stage_65;
  reg [31:0] dark_weights_update_0_stage_66;
  reg [31:0] dark_weights_update_0_stage_67;
  reg [31:0] dark_weights_update_0_stage_68;
  reg [31:0] dark_weights_update_0_stage_69;
  reg [31:0] dark_weights_update_0_stage_70;
  reg [31:0] dark_weights_update_0_stage_71;
  reg [31:0] dark_weights_update_0_stage_72;
  reg [31:0] dark_weights_update_0_stage_73;
  reg [31:0] dark_weights_update_0_stage_74;
  reg [31:0] dark_weights_update_0_stage_75;
  reg [31:0] dark_weights_update_0_stage_76;
  reg [31:0] dark_weights_update_0_stage_77;
  reg [31:0] dark_weights_update_0_stage_78;
  reg [31:0] dark_weights_update_0_stage_79;
  reg [31:0] dark_weights_update_0_stage_80;
  reg [31:0] dark_weights_update_0_stage_81;
  reg [31:0] dark_weights_update_0_stage_82;
  reg [31:0] dark_weights_update_0_stage_83;
  reg [31:0] dark_weights_update_0_stage_84;
  reg [31:0] dark_weights_update_0_stage_85;
  reg [31:0] dark_weights_update_0_stage_86;
  reg [31:0] dark_weights_update_0_stage_87;
  reg [31:0] dark_weights_update_0_stage_88;
  reg [31:0] dark_weights_update_0_stage_89;
  reg [31:0] dark_weights_update_0_stage_90;
  reg [31:0] dark_weights_update_0_stage_91;
  reg [31:0] dark_weights_update_0_stage_92;
  reg [31:0] dark_weights_update_0_stage_93;
  reg [31:0] dark_weights_update_0_stage_94;
  reg [31:0] dark_weights_update_0_stage_95;
  reg [31:0] dark_weights_update_0_stage_96;
  reg [31:0] dark_weights_update_0_stage_97;
  reg [31:0] dark_weights_update_0_stage_98;
  reg [31:0] dark_weights_update_0_stage_99;
  reg [31:0] dark_weights_update_0_stage_100;
  reg [31:0] dark_weights_update_0_stage_101;
  reg [31:0] dark_weights_update_0_stage_102;
  reg [31:0] dark_weights_update_0_stage_103;
  reg [31:0] dark_weights_update_0_stage_104;
  reg [31:0] dark_weights_update_0_stage_105;
  reg [31:0] dark_weights_update_0_stage_106;
  reg [31:0] dark_weights_update_0_stage_107;
  reg [31:0] dark_weights_update_0_stage_108;
  reg [31:0] dark_weights_update_0_stage_109;
  reg [31:0] dark_weights_update_0_stage_110;
  reg [31:0] dark_weights_update_0_stage_111;
  reg [31:0] dark_weights_update_0_stage_112;
  reg [31:0] dark_weights_update_0_stage_113;
  reg [31:0] dark_weights_update_0_stage_114;
  reg [31:0] dark_weights_update_0_stage_115;
  reg [31:0] dark_weights_update_0_stage_116;
  reg [31:0] dark_weights_update_0_stage_117;
  reg [31:0] dark_weights_update_0_stage_118;
  reg [31:0] dark_weights_update_0_stage_119;
  reg [31:0] dark_weights_update_0_stage_120;
  reg [31:0] dark_weights_update_0_stage_121;
  reg [31:0] dark_weights_update_0_stage_122;
  reg [31:0] dark_weights_update_0_stage_123;
  reg [31:0] dark_weights_update_0_stage_124;
  reg [31:0] dark_weights_update_0_stage_125;
  reg [31:0] dark_weights_update_0_stage_126;
  reg [31:0] dark_weights_update_0_stage_127;
  reg [31:0] dark_weights_update_0_stage_128;
  reg [31:0] dark_weights_update_0_stage_129;
  reg [31:0] dark_weights_update_0_stage_130;
  reg [31:0] dark_weights_update_0_stage_131;
  reg [31:0] dark_weights_update_0_stage_132;
  reg [31:0] dark_weights_update_0_stage_133;
  reg [31:0] dark_weights_update_0_stage_134;
  reg [31:0] dark_weights_update_0_stage_135;
  reg [31:0] dark_weights_update_0_stage_136;
  reg [31:0] dark_weights_update_0_stage_137;
  reg [31:0] dark_weights_update_0_stage_138;
  reg [31:0] dark_weights_update_0_stage_139;
  reg [31:0] dark_weights_update_0_stage_140;
  reg [31:0] dark_weights_update_0_stage_141;
  reg [31:0] dark_weights_update_0_stage_142;
  reg [31:0] dark_weights_update_0_stage_143;
  reg [31:0] dark_weights_update_0_stage_144;
  reg [31:0] dark_weights_update_0_stage_145;
  reg [31:0] dark_weights_update_0_stage_146;
  reg [31:0] dark_weights_update_0_stage_147;
  reg [31:0] dark_weights_update_0_stage_148;
  reg [31:0] dark_weights_update_0_stage_149;
  reg [31:0] dark_weights_update_0_stage_150;
  reg [31:0] dark_weights_update_0_stage_151;
  reg [31:0] dark_weights_update_0_stage_152;
  reg [31:0] dark_weights_update_0_stage_153;
  reg [31:0] dark_weights_update_0_stage_154;
  reg [31:0] dark_weights_update_0_stage_155;
  reg [31:0] dark_weights_update_0_stage_156;
  reg [31:0] dark_weights_update_0_stage_157;
  reg [31:0] dark_weights_update_0_stage_158;
  reg [31:0] dark_weights_update_0_stage_159;
  reg [31:0] dark_weights_update_0_stage_160;
  reg [31:0] dark_weights_update_0_stage_161;
  reg [31:0] dark_weights_update_0_stage_162;
  reg [31:0] dark_weights_update_0_stage_163;
  reg [31:0] dark_weights_update_0_stage_164;
  reg [31:0] dark_weights_update_0_stage_165;
  reg [31:0] dark_weights_update_0_stage_166;
  reg [31:0] dark_weights_update_0_stage_167;
  reg [31:0] dark_weights_update_0_stage_168;
  reg [31:0] dark_weights_update_0_stage_169;
  reg [31:0] dark_weights_update_0_stage_170;
  reg [31:0] dark_weights_update_0_stage_171;
  reg [31:0] dark_weights_update_0_stage_172;
  reg [31:0] dark_weights_update_0_stage_173;
  reg [31:0] dark_weights_update_0_stage_174;
  reg [31:0] dark_weights_update_0_stage_175;
  reg [31:0] dark_weights_update_0_stage_176;
  reg [31:0] dark_weights_update_0_stage_177;
  reg [31:0] dark_weights_update_0_stage_178;
  reg [31:0] dark_weights_update_0_stage_179;
  reg [31:0] dark_weights_update_0_stage_180;
  reg [31:0] dark_weights_update_0_stage_181;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_16;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_17;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_18;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_19;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_20;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_21;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_22;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_23;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_24;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_25;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_26;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_27;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_28;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_29;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_30;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_31;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_32;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_33;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_34;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_35;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_36;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_37;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_38;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_39;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_40;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_41;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_42;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_43;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_44;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_45;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_46;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_47;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_48;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_49;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_50;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_51;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_52;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_53;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_54;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_55;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_56;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_57;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_58;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_59;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_60;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_61;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_62;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_63;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_64;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_65;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_66;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_67;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_68;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_69;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_70;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_71;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_72;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_73;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_74;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_75;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_76;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_77;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_78;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_79;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_80;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_81;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_82;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_83;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_84;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_85;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_86;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_87;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_88;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_89;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_90;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_91;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_92;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_93;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_94;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_95;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_96;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_97;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_98;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_99;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_100;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_101;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_102;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_103;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_104;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_105;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_106;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_107;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_108;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_109;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_110;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_111;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_112;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_113;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_114;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_115;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_116;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_117;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_118;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_119;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_120;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_121;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_122;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_123;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_124;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_125;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_126;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_127;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_128;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_129;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_130;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_131;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_132;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_133;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_134;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_135;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_136;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_137;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_138;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_139;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_140;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_141;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_142;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_143;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_144;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_145;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_146;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_147;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_148;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_149;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_150;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_151;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_152;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_153;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_154;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_155;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_156;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_157;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_158;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_159;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_160;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_161;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_162;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_163;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_164;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_165;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_166;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_167;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_168;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_169;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_170;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_171;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_172;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_173;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_174;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_175;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_176;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_177;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_178;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_179;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_180;
  reg [31:0] dark_weights_dark_weights_update_0_write_write_9_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_86;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_87;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_88;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_89;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_90;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_91;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_92;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_93;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_2_update_0_stage_181;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_171;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_172;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_173;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_174;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_175;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_176;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_177;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_178;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_179;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_180;
  reg [31:0] final_merged_2_final_merged_1_update_0_read_read_120_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_87;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_88;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_89;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_90;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_91;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_92;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_93;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_181;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_172;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_173;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_174;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_175;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_176;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_177;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_178;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_179;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_180;
  reg [31:0] fused_level_1_final_merged_1_update_0_read_read_121_stage_181;
  reg [31:0] final_merged_1_update_0_stage_173;
  reg [31:0] final_merged_1_update_0_stage_174;
  reg [31:0] final_merged_1_update_0_stage_175;
  reg [31:0] final_merged_1_update_0_stage_176;
  reg [31:0] final_merged_1_update_0_stage_177;
  reg [31:0] final_merged_1_update_0_stage_178;
  reg [31:0] final_merged_1_update_0_stage_179;
  reg [31:0] final_merged_1_update_0_stage_180;
  reg [31:0] final_merged_1_update_0_stage_181;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_174;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_175;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_176;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_177;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_178;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_179;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_180;
  reg [31:0] final_merged_1_final_merged_1_update_0_write_write_122_stage_181;
  reg [31:0] in_in_update_0_write_write_1_stage_4;
  reg [31:0] in_in_update_0_write_write_1_stage_5;
  reg [31:0] in_in_update_0_write_write_1_stage_6;
  reg [31:0] in_in_update_0_write_write_1_stage_7;
  reg [31:0] in_in_update_0_write_write_1_stage_8;
  reg [31:0] in_in_update_0_write_write_1_stage_9;
  reg [31:0] in_in_update_0_write_write_1_stage_10;
  reg [31:0] in_in_update_0_write_write_1_stage_11;
  reg [31:0] in_in_update_0_write_write_1_stage_12;
  reg [31:0] in_in_update_0_write_write_1_stage_13;
  reg [31:0] in_in_update_0_write_write_1_stage_14;
  reg [31:0] in_in_update_0_write_write_1_stage_15;
  reg [31:0] in_in_update_0_write_write_1_stage_16;
  reg [31:0] in_in_update_0_write_write_1_stage_17;
  reg [31:0] in_in_update_0_write_write_1_stage_18;
  reg [31:0] in_in_update_0_write_write_1_stage_19;
  reg [31:0] in_in_update_0_write_write_1_stage_20;
  reg [31:0] in_in_update_0_write_write_1_stage_21;
  reg [31:0] in_in_update_0_write_write_1_stage_22;
  reg [31:0] in_in_update_0_write_write_1_stage_23;
  reg [31:0] in_in_update_0_write_write_1_stage_24;
  reg [31:0] in_in_update_0_write_write_1_stage_25;
  reg [31:0] in_in_update_0_write_write_1_stage_26;
  reg [31:0] in_in_update_0_write_write_1_stage_27;
  reg [31:0] in_in_update_0_write_write_1_stage_28;
  reg [31:0] in_in_update_0_write_write_1_stage_29;
  reg [31:0] in_in_update_0_write_write_1_stage_30;
  reg [31:0] in_in_update_0_write_write_1_stage_31;
  reg [31:0] in_in_update_0_write_write_1_stage_32;
  reg [31:0] in_in_update_0_write_write_1_stage_33;
  reg [31:0] in_in_update_0_write_write_1_stage_34;
  reg [31:0] in_in_update_0_write_write_1_stage_35;
  reg [31:0] in_in_update_0_write_write_1_stage_36;
  reg [31:0] in_in_update_0_write_write_1_stage_37;
  reg [31:0] in_in_update_0_write_write_1_stage_38;
  reg [31:0] in_in_update_0_write_write_1_stage_39;
  reg [31:0] in_in_update_0_write_write_1_stage_40;
  reg [31:0] in_in_update_0_write_write_1_stage_41;
  reg [31:0] in_in_update_0_write_write_1_stage_42;
  reg [31:0] in_in_update_0_write_write_1_stage_43;
  reg [31:0] in_in_update_0_write_write_1_stage_44;
  reg [31:0] in_in_update_0_write_write_1_stage_45;
  reg [31:0] in_in_update_0_write_write_1_stage_46;
  reg [31:0] in_in_update_0_write_write_1_stage_47;
  reg [31:0] in_in_update_0_write_write_1_stage_48;
  reg [31:0] in_in_update_0_write_write_1_stage_49;
  reg [31:0] in_in_update_0_write_write_1_stage_50;
  reg [31:0] in_in_update_0_write_write_1_stage_51;
  reg [31:0] in_in_update_0_write_write_1_stage_52;
  reg [31:0] in_in_update_0_write_write_1_stage_53;
  reg [31:0] in_in_update_0_write_write_1_stage_54;
  reg [31:0] in_in_update_0_write_write_1_stage_55;
  reg [31:0] in_in_update_0_write_write_1_stage_56;
  reg [31:0] in_in_update_0_write_write_1_stage_57;
  reg [31:0] in_in_update_0_write_write_1_stage_58;
  reg [31:0] in_in_update_0_write_write_1_stage_59;
  reg [31:0] in_in_update_0_write_write_1_stage_60;
  reg [31:0] in_in_update_0_write_write_1_stage_61;
  reg [31:0] in_in_update_0_write_write_1_stage_62;
  reg [31:0] in_in_update_0_write_write_1_stage_63;
  reg [31:0] in_in_update_0_write_write_1_stage_64;
  reg [31:0] in_in_update_0_write_write_1_stage_65;
  reg [31:0] in_in_update_0_write_write_1_stage_66;
  reg [31:0] in_in_update_0_write_write_1_stage_67;
  reg [31:0] in_in_update_0_write_write_1_stage_68;
  reg [31:0] in_in_update_0_write_write_1_stage_69;
  reg [31:0] in_in_update_0_write_write_1_stage_70;
  reg [31:0] in_in_update_0_write_write_1_stage_71;
  reg [31:0] in_in_update_0_write_write_1_stage_72;
  reg [31:0] in_in_update_0_write_write_1_stage_73;
  reg [31:0] in_in_update_0_write_write_1_stage_74;
  reg [31:0] in_in_update_0_write_write_1_stage_75;
  reg [31:0] in_in_update_0_write_write_1_stage_76;
  reg [31:0] in_in_update_0_write_write_1_stage_77;
  reg [31:0] in_in_update_0_write_write_1_stage_78;
  reg [31:0] in_in_update_0_write_write_1_stage_79;
  reg [31:0] in_in_update_0_write_write_1_stage_80;
  reg [31:0] in_in_update_0_write_write_1_stage_81;
  reg [31:0] in_in_update_0_write_write_1_stage_82;
  reg [31:0] in_in_update_0_write_write_1_stage_83;
  reg [31:0] in_in_update_0_write_write_1_stage_84;
  reg [31:0] in_in_update_0_write_write_1_stage_85;
  reg [31:0] in_in_update_0_write_write_1_stage_86;
  reg [31:0] in_in_update_0_write_write_1_stage_87;
  reg [31:0] in_in_update_0_write_write_1_stage_88;
  reg [31:0] in_in_update_0_write_write_1_stage_89;
  reg [31:0] in_in_update_0_write_write_1_stage_90;
  reg [31:0] in_in_update_0_write_write_1_stage_91;
  reg [31:0] in_in_update_0_write_write_1_stage_92;
  reg [31:0] in_in_update_0_write_write_1_stage_93;
  reg [31:0] in_in_update_0_write_write_1_stage_94;
  reg [31:0] in_in_update_0_write_write_1_stage_95;
  reg [31:0] in_in_update_0_write_write_1_stage_96;
  reg [31:0] in_in_update_0_write_write_1_stage_97;
  reg [31:0] in_in_update_0_write_write_1_stage_98;
  reg [31:0] in_in_update_0_write_write_1_stage_99;
  reg [31:0] in_in_update_0_write_write_1_stage_100;
  reg [31:0] in_in_update_0_write_write_1_stage_101;
  reg [31:0] in_in_update_0_write_write_1_stage_102;
  reg [31:0] in_in_update_0_write_write_1_stage_103;
  reg [31:0] in_in_update_0_write_write_1_stage_104;
  reg [31:0] in_in_update_0_write_write_1_stage_105;
  reg [31:0] in_in_update_0_write_write_1_stage_106;
  reg [31:0] in_in_update_0_write_write_1_stage_107;
  reg [31:0] in_in_update_0_write_write_1_stage_108;
  reg [31:0] in_in_update_0_write_write_1_stage_109;
  reg [31:0] in_in_update_0_write_write_1_stage_110;
  reg [31:0] in_in_update_0_write_write_1_stage_111;
  reg [31:0] in_in_update_0_write_write_1_stage_112;
  reg [31:0] in_in_update_0_write_write_1_stage_113;
  reg [31:0] in_in_update_0_write_write_1_stage_114;
  reg [31:0] in_in_update_0_write_write_1_stage_115;
  reg [31:0] in_in_update_0_write_write_1_stage_116;
  reg [31:0] in_in_update_0_write_write_1_stage_117;
  reg [31:0] in_in_update_0_write_write_1_stage_118;
  reg [31:0] in_in_update_0_write_write_1_stage_119;
  reg [31:0] in_in_update_0_write_write_1_stage_120;
  reg [31:0] in_in_update_0_write_write_1_stage_121;
  reg [31:0] in_in_update_0_write_write_1_stage_122;
  reg [31:0] in_in_update_0_write_write_1_stage_123;
  reg [31:0] in_in_update_0_write_write_1_stage_124;
  reg [31:0] in_in_update_0_write_write_1_stage_125;
  reg [31:0] in_in_update_0_write_write_1_stage_126;
  reg [31:0] in_in_update_0_write_write_1_stage_127;
  reg [31:0] in_in_update_0_write_write_1_stage_128;
  reg [31:0] in_in_update_0_write_write_1_stage_129;
  reg [31:0] in_in_update_0_write_write_1_stage_130;
  reg [31:0] in_in_update_0_write_write_1_stage_131;
  reg [31:0] in_in_update_0_write_write_1_stage_132;
  reg [31:0] in_in_update_0_write_write_1_stage_133;
  reg [31:0] in_in_update_0_write_write_1_stage_134;
  reg [31:0] in_in_update_0_write_write_1_stage_135;
  reg [31:0] in_in_update_0_write_write_1_stage_136;
  reg [31:0] in_in_update_0_write_write_1_stage_137;
  reg [31:0] in_in_update_0_write_write_1_stage_138;
  reg [31:0] in_in_update_0_write_write_1_stage_139;
  reg [31:0] in_in_update_0_write_write_1_stage_140;
  reg [31:0] in_in_update_0_write_write_1_stage_141;
  reg [31:0] in_in_update_0_write_write_1_stage_142;
  reg [31:0] in_in_update_0_write_write_1_stage_143;
  reg [31:0] in_in_update_0_write_write_1_stage_144;
  reg [31:0] in_in_update_0_write_write_1_stage_145;
  reg [31:0] in_in_update_0_write_write_1_stage_146;
  reg [31:0] in_in_update_0_write_write_1_stage_147;
  reg [31:0] in_in_update_0_write_write_1_stage_148;
  reg [31:0] in_in_update_0_write_write_1_stage_149;
  reg [31:0] in_in_update_0_write_write_1_stage_150;
  reg [31:0] in_in_update_0_write_write_1_stage_151;
  reg [31:0] in_in_update_0_write_write_1_stage_152;
  reg [31:0] in_in_update_0_write_write_1_stage_153;
  reg [31:0] in_in_update_0_write_write_1_stage_154;
  reg [31:0] in_in_update_0_write_write_1_stage_155;
  reg [31:0] in_in_update_0_write_write_1_stage_156;
  reg [31:0] in_in_update_0_write_write_1_stage_157;
  reg [31:0] in_in_update_0_write_write_1_stage_158;
  reg [31:0] in_in_update_0_write_write_1_stage_159;
  reg [31:0] in_in_update_0_write_write_1_stage_160;
  reg [31:0] in_in_update_0_write_write_1_stage_161;
  reg [31:0] in_in_update_0_write_write_1_stage_162;
  reg [31:0] in_in_update_0_write_write_1_stage_163;
  reg [31:0] in_in_update_0_write_write_1_stage_164;
  reg [31:0] in_in_update_0_write_write_1_stage_165;
  reg [31:0] in_in_update_0_write_write_1_stage_166;
  reg [31:0] in_in_update_0_write_write_1_stage_167;
  reg [31:0] in_in_update_0_write_write_1_stage_168;
  reg [31:0] in_in_update_0_write_write_1_stage_169;
  reg [31:0] in_in_update_0_write_write_1_stage_170;
  reg [31:0] in_in_update_0_write_write_1_stage_171;
  reg [31:0] in_in_update_0_write_write_1_stage_172;
  reg [31:0] in_in_update_0_write_write_1_stage_173;
  reg [31:0] in_in_update_0_write_write_1_stage_174;
  reg [31:0] in_in_update_0_write_write_1_stage_175;
  reg [31:0] in_in_update_0_write_write_1_stage_176;
  reg [31:0] in_in_update_0_write_write_1_stage_177;
  reg [31:0] in_in_update_0_write_write_1_stage_178;
  reg [31:0] in_in_update_0_write_write_1_stage_179;
  reg [31:0] in_in_update_0_write_write_1_stage_180;
  reg [31:0] in_in_update_0_write_write_1_stage_181;
  reg [31:0] in_bright_update_0_read_read_2_stage_5;
  reg [31:0] in_bright_update_0_read_read_2_stage_6;
  reg [31:0] in_bright_update_0_read_read_2_stage_7;
  reg [31:0] in_bright_update_0_read_read_2_stage_8;
  reg [31:0] in_bright_update_0_read_read_2_stage_9;
  reg [31:0] in_bright_update_0_read_read_2_stage_10;
  reg [31:0] in_bright_update_0_read_read_2_stage_11;
  reg [31:0] in_bright_update_0_read_read_2_stage_12;
  reg [31:0] in_bright_update_0_read_read_2_stage_13;
  reg [31:0] in_bright_update_0_read_read_2_stage_14;
  reg [31:0] in_bright_update_0_read_read_2_stage_15;
  reg [31:0] in_bright_update_0_read_read_2_stage_16;
  reg [31:0] in_bright_update_0_read_read_2_stage_17;
  reg [31:0] in_bright_update_0_read_read_2_stage_18;
  reg [31:0] in_bright_update_0_read_read_2_stage_19;
  reg [31:0] in_bright_update_0_read_read_2_stage_20;
  reg [31:0] in_bright_update_0_read_read_2_stage_21;
  reg [31:0] in_bright_update_0_read_read_2_stage_22;
  reg [31:0] in_bright_update_0_read_read_2_stage_23;
  reg [31:0] in_bright_update_0_read_read_2_stage_24;
  reg [31:0] in_bright_update_0_read_read_2_stage_25;
  reg [31:0] in_bright_update_0_read_read_2_stage_26;
  reg [31:0] in_bright_update_0_read_read_2_stage_27;
  reg [31:0] in_bright_update_0_read_read_2_stage_28;
  reg [31:0] in_bright_update_0_read_read_2_stage_29;
  reg [31:0] in_bright_update_0_read_read_2_stage_30;
  reg [31:0] in_bright_update_0_read_read_2_stage_31;
  reg [31:0] in_bright_update_0_read_read_2_stage_32;
  reg [31:0] in_bright_update_0_read_read_2_stage_33;
  reg [31:0] in_bright_update_0_read_read_2_stage_34;
  reg [31:0] in_bright_update_0_read_read_2_stage_35;
  reg [31:0] in_bright_update_0_read_read_2_stage_36;
  reg [31:0] in_bright_update_0_read_read_2_stage_37;
  reg [31:0] in_bright_update_0_read_read_2_stage_38;
  reg [31:0] in_bright_update_0_read_read_2_stage_39;
  reg [31:0] in_bright_update_0_read_read_2_stage_40;
  reg [31:0] in_bright_update_0_read_read_2_stage_41;
  reg [31:0] in_bright_update_0_read_read_2_stage_42;
  reg [31:0] in_bright_update_0_read_read_2_stage_43;
  reg [31:0] in_bright_update_0_read_read_2_stage_44;
  reg [31:0] in_bright_update_0_read_read_2_stage_45;
  reg [31:0] in_bright_update_0_read_read_2_stage_46;
  reg [31:0] in_bright_update_0_read_read_2_stage_47;
  reg [31:0] in_bright_update_0_read_read_2_stage_48;
  reg [31:0] in_bright_update_0_read_read_2_stage_49;
  reg [31:0] in_bright_update_0_read_read_2_stage_50;
  reg [31:0] in_bright_update_0_read_read_2_stage_51;
  reg [31:0] in_bright_update_0_read_read_2_stage_52;
  reg [31:0] in_bright_update_0_read_read_2_stage_53;
  reg [31:0] in_bright_update_0_read_read_2_stage_54;
  reg [31:0] in_bright_update_0_read_read_2_stage_55;
  reg [31:0] in_bright_update_0_read_read_2_stage_56;
  reg [31:0] in_bright_update_0_read_read_2_stage_57;
  reg [31:0] in_bright_update_0_read_read_2_stage_58;
  reg [31:0] in_bright_update_0_read_read_2_stage_59;
  reg [31:0] in_bright_update_0_read_read_2_stage_60;
  reg [31:0] in_bright_update_0_read_read_2_stage_61;
  reg [31:0] in_bright_update_0_read_read_2_stage_62;
  reg [31:0] in_bright_update_0_read_read_2_stage_63;
  reg [31:0] in_bright_update_0_read_read_2_stage_64;
  reg [31:0] in_bright_update_0_read_read_2_stage_65;
  reg [31:0] in_bright_update_0_read_read_2_stage_66;
  reg [31:0] in_bright_update_0_read_read_2_stage_67;
  reg [31:0] in_bright_update_0_read_read_2_stage_68;
  reg [31:0] in_bright_update_0_read_read_2_stage_69;
  reg [31:0] in_bright_update_0_read_read_2_stage_70;
  reg [31:0] in_bright_update_0_read_read_2_stage_71;
  reg [31:0] in_bright_update_0_read_read_2_stage_72;
  reg [31:0] in_bright_update_0_read_read_2_stage_73;
  reg [31:0] in_bright_update_0_read_read_2_stage_74;
  reg [31:0] in_bright_update_0_read_read_2_stage_75;
  reg [31:0] in_bright_update_0_read_read_2_stage_76;
  reg [31:0] in_bright_update_0_read_read_2_stage_77;
  reg [31:0] in_bright_update_0_read_read_2_stage_78;
  reg [31:0] in_bright_update_0_read_read_2_stage_79;
  reg [31:0] in_bright_update_0_read_read_2_stage_80;
  reg [31:0] in_bright_update_0_read_read_2_stage_81;
  reg [31:0] in_bright_update_0_read_read_2_stage_82;
  reg [31:0] in_bright_update_0_read_read_2_stage_83;
  reg [31:0] in_bright_update_0_read_read_2_stage_84;
  reg [31:0] in_bright_update_0_read_read_2_stage_85;
  reg [31:0] in_bright_update_0_read_read_2_stage_86;
  reg [31:0] in_bright_update_0_read_read_2_stage_87;
  reg [31:0] in_bright_update_0_read_read_2_stage_88;
  reg [31:0] in_bright_update_0_read_read_2_stage_89;
  reg [31:0] in_bright_update_0_read_read_2_stage_90;
  reg [31:0] in_bright_update_0_read_read_2_stage_91;
  reg [31:0] in_bright_update_0_read_read_2_stage_92;
  reg [31:0] in_bright_update_0_read_read_2_stage_93;
  reg [31:0] in_bright_update_0_read_read_2_stage_94;
  reg [31:0] in_bright_update_0_read_read_2_stage_95;
  reg [31:0] in_bright_update_0_read_read_2_stage_96;
  reg [31:0] in_bright_update_0_read_read_2_stage_97;
  reg [31:0] in_bright_update_0_read_read_2_stage_98;
  reg [31:0] in_bright_update_0_read_read_2_stage_99;
  reg [31:0] in_bright_update_0_read_read_2_stage_100;
  reg [31:0] in_bright_update_0_read_read_2_stage_101;
  reg [31:0] in_bright_update_0_read_read_2_stage_102;
  reg [31:0] in_bright_update_0_read_read_2_stage_103;
  reg [31:0] in_bright_update_0_read_read_2_stage_104;
  reg [31:0] in_bright_update_0_read_read_2_stage_105;
  reg [31:0] in_bright_update_0_read_read_2_stage_106;
  reg [31:0] in_bright_update_0_read_read_2_stage_107;
  reg [31:0] in_bright_update_0_read_read_2_stage_108;
  reg [31:0] in_bright_update_0_read_read_2_stage_109;
  reg [31:0] in_bright_update_0_read_read_2_stage_110;
  reg [31:0] in_bright_update_0_read_read_2_stage_111;
  reg [31:0] in_bright_update_0_read_read_2_stage_112;
  reg [31:0] in_bright_update_0_read_read_2_stage_113;
  reg [31:0] in_bright_update_0_read_read_2_stage_114;
  reg [31:0] in_bright_update_0_read_read_2_stage_115;
  reg [31:0] in_bright_update_0_read_read_2_stage_116;
  reg [31:0] in_bright_update_0_read_read_2_stage_117;
  reg [31:0] in_bright_update_0_read_read_2_stage_118;
  reg [31:0] in_bright_update_0_read_read_2_stage_119;
  reg [31:0] in_bright_update_0_read_read_2_stage_120;
  reg [31:0] in_bright_update_0_read_read_2_stage_121;
  reg [31:0] in_bright_update_0_read_read_2_stage_122;
  reg [31:0] in_bright_update_0_read_read_2_stage_123;
  reg [31:0] in_bright_update_0_read_read_2_stage_124;
  reg [31:0] in_bright_update_0_read_read_2_stage_125;
  reg [31:0] in_bright_update_0_read_read_2_stage_126;
  reg [31:0] in_bright_update_0_read_read_2_stage_127;
  reg [31:0] in_bright_update_0_read_read_2_stage_128;
  reg [31:0] in_bright_update_0_read_read_2_stage_129;
  reg [31:0] in_bright_update_0_read_read_2_stage_130;
  reg [31:0] in_bright_update_0_read_read_2_stage_131;
  reg [31:0] in_bright_update_0_read_read_2_stage_132;
  reg [31:0] in_bright_update_0_read_read_2_stage_133;
  reg [31:0] in_bright_update_0_read_read_2_stage_134;
  reg [31:0] in_bright_update_0_read_read_2_stage_135;
  reg [31:0] in_bright_update_0_read_read_2_stage_136;
  reg [31:0] in_bright_update_0_read_read_2_stage_137;
  reg [31:0] in_bright_update_0_read_read_2_stage_138;
  reg [31:0] in_bright_update_0_read_read_2_stage_139;
  reg [31:0] in_bright_update_0_read_read_2_stage_140;
  reg [31:0] in_bright_update_0_read_read_2_stage_141;
  reg [31:0] in_bright_update_0_read_read_2_stage_142;
  reg [31:0] in_bright_update_0_read_read_2_stage_143;
  reg [31:0] in_bright_update_0_read_read_2_stage_144;
  reg [31:0] in_bright_update_0_read_read_2_stage_145;
  reg [31:0] in_bright_update_0_read_read_2_stage_146;
  reg [31:0] in_bright_update_0_read_read_2_stage_147;
  reg [31:0] in_bright_update_0_read_read_2_stage_148;
  reg [31:0] in_bright_update_0_read_read_2_stage_149;
  reg [31:0] in_bright_update_0_read_read_2_stage_150;
  reg [31:0] in_bright_update_0_read_read_2_stage_151;
  reg [31:0] in_bright_update_0_read_read_2_stage_152;
  reg [31:0] in_bright_update_0_read_read_2_stage_153;
  reg [31:0] in_bright_update_0_read_read_2_stage_154;
  reg [31:0] in_bright_update_0_read_read_2_stage_155;
  reg [31:0] in_bright_update_0_read_read_2_stage_156;
  reg [31:0] in_bright_update_0_read_read_2_stage_157;
  reg [31:0] in_bright_update_0_read_read_2_stage_158;
  reg [31:0] in_bright_update_0_read_read_2_stage_159;
  reg [31:0] in_bright_update_0_read_read_2_stage_160;
  reg [31:0] in_bright_update_0_read_read_2_stage_161;
  reg [31:0] in_bright_update_0_read_read_2_stage_162;
  reg [31:0] in_bright_update_0_read_read_2_stage_163;
  reg [31:0] in_bright_update_0_read_read_2_stage_164;
  reg [31:0] in_bright_update_0_read_read_2_stage_165;
  reg [31:0] in_bright_update_0_read_read_2_stage_166;
  reg [31:0] in_bright_update_0_read_read_2_stage_167;
  reg [31:0] in_bright_update_0_read_read_2_stage_168;
  reg [31:0] in_bright_update_0_read_read_2_stage_169;
  reg [31:0] in_bright_update_0_read_read_2_stage_170;
  reg [31:0] in_bright_update_0_read_read_2_stage_171;
  reg [31:0] in_bright_update_0_read_read_2_stage_172;
  reg [31:0] in_bright_update_0_read_read_2_stage_173;
  reg [31:0] in_bright_update_0_read_read_2_stage_174;
  reg [31:0] in_bright_update_0_read_read_2_stage_175;
  reg [31:0] in_bright_update_0_read_read_2_stage_176;
  reg [31:0] in_bright_update_0_read_read_2_stage_177;
  reg [31:0] in_bright_update_0_read_read_2_stage_178;
  reg [31:0] in_bright_update_0_read_read_2_stage_179;
  reg [31:0] in_bright_update_0_read_read_2_stage_180;
  reg [31:0] in_bright_update_0_read_read_2_stage_181;
  reg [31:0] bright_update_0_stage_6;
  reg [31:0] bright_update_0_stage_7;
  reg [31:0] bright_update_0_stage_8;
  reg [31:0] bright_update_0_stage_9;
  reg [31:0] bright_update_0_stage_10;
  reg [31:0] bright_update_0_stage_11;
  reg [31:0] bright_update_0_stage_12;
  reg [31:0] bright_update_0_stage_13;
  reg [31:0] bright_update_0_stage_14;
  reg [31:0] bright_update_0_stage_15;
  reg [31:0] bright_update_0_stage_16;
  reg [31:0] bright_update_0_stage_17;
  reg [31:0] bright_update_0_stage_18;
  reg [31:0] bright_update_0_stage_19;
  reg [31:0] bright_update_0_stage_20;
  reg [31:0] bright_update_0_stage_21;
  reg [31:0] bright_update_0_stage_22;
  reg [31:0] bright_update_0_stage_23;
  reg [31:0] bright_update_0_stage_24;
  reg [31:0] bright_update_0_stage_25;
  reg [31:0] bright_update_0_stage_26;
  reg [31:0] bright_update_0_stage_27;
  reg [31:0] bright_update_0_stage_28;
  reg [31:0] bright_update_0_stage_29;
  reg [31:0] bright_update_0_stage_30;
  reg [31:0] bright_update_0_stage_31;
  reg [31:0] bright_update_0_stage_32;
  reg [31:0] bright_update_0_stage_33;
  reg [31:0] bright_update_0_stage_34;
  reg [31:0] bright_update_0_stage_35;
  reg [31:0] bright_update_0_stage_36;
  reg [31:0] bright_update_0_stage_37;
  reg [31:0] bright_update_0_stage_38;
  reg [31:0] bright_update_0_stage_39;
  reg [31:0] bright_update_0_stage_40;
  reg [31:0] bright_update_0_stage_41;
  reg [31:0] bright_update_0_stage_42;
  reg [31:0] bright_update_0_stage_43;
  reg [31:0] bright_update_0_stage_44;
  reg [31:0] bright_update_0_stage_45;
  reg [31:0] bright_update_0_stage_46;
  reg [31:0] bright_update_0_stage_47;
  reg [31:0] bright_update_0_stage_48;
  reg [31:0] bright_update_0_stage_49;
  reg [31:0] bright_update_0_stage_50;
  reg [31:0] bright_update_0_stage_51;
  reg [31:0] bright_update_0_stage_52;
  reg [31:0] bright_update_0_stage_53;
  reg [31:0] bright_update_0_stage_54;
  reg [31:0] bright_update_0_stage_55;
  reg [31:0] bright_update_0_stage_56;
  reg [31:0] bright_update_0_stage_57;
  reg [31:0] bright_update_0_stage_58;
  reg [31:0] bright_update_0_stage_59;
  reg [31:0] bright_update_0_stage_60;
  reg [31:0] bright_update_0_stage_61;
  reg [31:0] bright_update_0_stage_62;
  reg [31:0] bright_update_0_stage_63;
  reg [31:0] bright_update_0_stage_64;
  reg [31:0] bright_update_0_stage_65;
  reg [31:0] bright_update_0_stage_66;
  reg [31:0] bright_update_0_stage_67;
  reg [31:0] bright_update_0_stage_68;
  reg [31:0] bright_update_0_stage_69;
  reg [31:0] bright_update_0_stage_70;
  reg [31:0] bright_update_0_stage_71;
  reg [31:0] bright_update_0_stage_72;
  reg [31:0] bright_update_0_stage_73;
  reg [31:0] bright_update_0_stage_74;
  reg [31:0] bright_update_0_stage_75;
  reg [31:0] bright_update_0_stage_76;
  reg [31:0] bright_update_0_stage_77;
  reg [31:0] bright_update_0_stage_78;
  reg [31:0] bright_update_0_stage_79;
  reg [31:0] bright_update_0_stage_80;
  reg [31:0] bright_update_0_stage_81;
  reg [31:0] bright_update_0_stage_82;
  reg [31:0] bright_update_0_stage_83;
  reg [31:0] bright_update_0_stage_84;
  reg [31:0] bright_update_0_stage_85;
  reg [31:0] bright_update_0_stage_86;
  reg [31:0] bright_update_0_stage_87;
  reg [31:0] bright_update_0_stage_88;
  reg [31:0] bright_update_0_stage_89;
  reg [31:0] bright_update_0_stage_90;
  reg [31:0] bright_update_0_stage_91;
  reg [31:0] bright_update_0_stage_92;
  reg [31:0] bright_update_0_stage_93;
  reg [31:0] bright_update_0_stage_94;
  reg [31:0] bright_update_0_stage_95;
  reg [31:0] bright_update_0_stage_96;
  reg [31:0] bright_update_0_stage_97;
  reg [31:0] bright_update_0_stage_98;
  reg [31:0] bright_update_0_stage_99;
  reg [31:0] bright_update_0_stage_100;
  reg [31:0] bright_update_0_stage_101;
  reg [31:0] bright_update_0_stage_102;
  reg [31:0] bright_update_0_stage_103;
  reg [31:0] bright_update_0_stage_104;
  reg [31:0] bright_update_0_stage_105;
  reg [31:0] bright_update_0_stage_106;
  reg [31:0] bright_update_0_stage_107;
  reg [31:0] bright_update_0_stage_108;
  reg [31:0] bright_update_0_stage_109;
  reg [31:0] bright_update_0_stage_110;
  reg [31:0] bright_update_0_stage_111;
  reg [31:0] bright_update_0_stage_112;
  reg [31:0] bright_update_0_stage_113;
  reg [31:0] bright_update_0_stage_114;
  reg [31:0] bright_update_0_stage_115;
  reg [31:0] bright_update_0_stage_116;
  reg [31:0] bright_update_0_stage_117;
  reg [31:0] bright_update_0_stage_118;
  reg [31:0] bright_update_0_stage_119;
  reg [31:0] bright_update_0_stage_120;
  reg [31:0] bright_update_0_stage_121;
  reg [31:0] bright_update_0_stage_122;
  reg [31:0] bright_update_0_stage_123;
  reg [31:0] bright_update_0_stage_124;
  reg [31:0] bright_update_0_stage_125;
  reg [31:0] bright_update_0_stage_126;
  reg [31:0] bright_update_0_stage_127;
  reg [31:0] bright_update_0_stage_128;
  reg [31:0] bright_update_0_stage_129;
  reg [31:0] bright_update_0_stage_130;
  reg [31:0] bright_update_0_stage_131;
  reg [31:0] bright_update_0_stage_132;
  reg [31:0] bright_update_0_stage_133;
  reg [31:0] bright_update_0_stage_134;
  reg [31:0] bright_update_0_stage_135;
  reg [31:0] bright_update_0_stage_136;
  reg [31:0] bright_update_0_stage_137;
  reg [31:0] bright_update_0_stage_138;
  reg [31:0] bright_update_0_stage_139;
  reg [31:0] bright_update_0_stage_140;
  reg [31:0] bright_update_0_stage_141;
  reg [31:0] bright_update_0_stage_142;
  reg [31:0] bright_update_0_stage_143;
  reg [31:0] bright_update_0_stage_144;
  reg [31:0] bright_update_0_stage_145;
  reg [31:0] bright_update_0_stage_146;
  reg [31:0] bright_update_0_stage_147;
  reg [31:0] bright_update_0_stage_148;
  reg [31:0] bright_update_0_stage_149;
  reg [31:0] bright_update_0_stage_150;
  reg [31:0] bright_update_0_stage_151;
  reg [31:0] bright_update_0_stage_152;
  reg [31:0] bright_update_0_stage_153;
  reg [31:0] bright_update_0_stage_154;
  reg [31:0] bright_update_0_stage_155;
  reg [31:0] bright_update_0_stage_156;
  reg [31:0] bright_update_0_stage_157;
  reg [31:0] bright_update_0_stage_158;
  reg [31:0] bright_update_0_stage_159;
  reg [31:0] bright_update_0_stage_160;
  reg [31:0] bright_update_0_stage_161;
  reg [31:0] bright_update_0_stage_162;
  reg [31:0] bright_update_0_stage_163;
  reg [31:0] bright_update_0_stage_164;
  reg [31:0] bright_update_0_stage_165;
  reg [31:0] bright_update_0_stage_166;
  reg [31:0] bright_update_0_stage_167;
  reg [31:0] bright_update_0_stage_168;
  reg [31:0] bright_update_0_stage_169;
  reg [31:0] bright_update_0_stage_170;
  reg [31:0] bright_update_0_stage_171;
  reg [31:0] bright_update_0_stage_172;
  reg [31:0] bright_update_0_stage_173;
  reg [31:0] bright_update_0_stage_174;
  reg [31:0] bright_update_0_stage_175;
  reg [31:0] bright_update_0_stage_176;
  reg [31:0] bright_update_0_stage_177;
  reg [31:0] bright_update_0_stage_178;
  reg [31:0] bright_update_0_stage_179;
  reg [31:0] bright_update_0_stage_180;
  reg [31:0] bright_update_0_stage_181;
  reg [31:0] bright_bright_update_0_write_write_3_stage_7;
  reg [31:0] bright_bright_update_0_write_write_3_stage_8;
  reg [31:0] bright_bright_update_0_write_write_3_stage_9;
  reg [31:0] bright_bright_update_0_write_write_3_stage_10;
  reg [31:0] bright_bright_update_0_write_write_3_stage_11;
  reg [31:0] bright_bright_update_0_write_write_3_stage_12;
  reg [31:0] bright_bright_update_0_write_write_3_stage_13;
  reg [31:0] bright_bright_update_0_write_write_3_stage_14;
  reg [31:0] bright_bright_update_0_write_write_3_stage_15;
  reg [31:0] bright_bright_update_0_write_write_3_stage_16;
  reg [31:0] bright_bright_update_0_write_write_3_stage_17;
  reg [31:0] bright_bright_update_0_write_write_3_stage_18;
  reg [31:0] bright_bright_update_0_write_write_3_stage_19;
  reg [31:0] bright_bright_update_0_write_write_3_stage_20;
  reg [31:0] bright_bright_update_0_write_write_3_stage_21;
  reg [31:0] bright_bright_update_0_write_write_3_stage_22;
  reg [31:0] bright_bright_update_0_write_write_3_stage_23;
  reg [31:0] bright_bright_update_0_write_write_3_stage_24;
  reg [31:0] bright_bright_update_0_write_write_3_stage_25;
  reg [31:0] bright_bright_update_0_write_write_3_stage_26;
  reg [31:0] bright_bright_update_0_write_write_3_stage_27;
  reg [31:0] bright_bright_update_0_write_write_3_stage_28;
  reg [31:0] bright_bright_update_0_write_write_3_stage_29;
  reg [31:0] bright_bright_update_0_write_write_3_stage_30;
  reg [31:0] bright_bright_update_0_write_write_3_stage_31;
  reg [31:0] bright_bright_update_0_write_write_3_stage_32;
  reg [31:0] bright_bright_update_0_write_write_3_stage_33;
  reg [31:0] bright_bright_update_0_write_write_3_stage_34;
  reg [31:0] bright_bright_update_0_write_write_3_stage_35;
  reg [31:0] bright_bright_update_0_write_write_3_stage_36;
  reg [31:0] bright_bright_update_0_write_write_3_stage_37;
  reg [31:0] bright_bright_update_0_write_write_3_stage_38;
  reg [31:0] bright_bright_update_0_write_write_3_stage_39;
  reg [31:0] bright_bright_update_0_write_write_3_stage_40;
  reg [31:0] bright_bright_update_0_write_write_3_stage_41;
  reg [31:0] bright_bright_update_0_write_write_3_stage_42;
  reg [31:0] bright_bright_update_0_write_write_3_stage_43;
  reg [31:0] bright_bright_update_0_write_write_3_stage_44;
  reg [31:0] bright_bright_update_0_write_write_3_stage_45;
  reg [31:0] bright_bright_update_0_write_write_3_stage_46;
  reg [31:0] bright_bright_update_0_write_write_3_stage_47;
  reg [31:0] bright_bright_update_0_write_write_3_stage_48;
  reg [31:0] bright_bright_update_0_write_write_3_stage_49;
  reg [31:0] bright_bright_update_0_write_write_3_stage_50;
  reg [31:0] bright_bright_update_0_write_write_3_stage_51;
  reg [31:0] bright_bright_update_0_write_write_3_stage_52;
  reg [31:0] bright_bright_update_0_write_write_3_stage_53;
  reg [31:0] bright_bright_update_0_write_write_3_stage_54;
  reg [31:0] bright_bright_update_0_write_write_3_stage_55;
  reg [31:0] bright_bright_update_0_write_write_3_stage_56;
  reg [31:0] bright_bright_update_0_write_write_3_stage_57;
  reg [31:0] bright_bright_update_0_write_write_3_stage_58;
  reg [31:0] bright_bright_update_0_write_write_3_stage_59;
  reg [31:0] bright_bright_update_0_write_write_3_stage_60;
  reg [31:0] bright_bright_update_0_write_write_3_stage_61;
  reg [31:0] bright_bright_update_0_write_write_3_stage_62;
  reg [31:0] bright_bright_update_0_write_write_3_stage_63;
  reg [31:0] bright_bright_update_0_write_write_3_stage_64;
  reg [31:0] bright_bright_update_0_write_write_3_stage_65;
  reg [31:0] bright_bright_update_0_write_write_3_stage_66;
  reg [31:0] bright_bright_update_0_write_write_3_stage_67;
  reg [31:0] bright_bright_update_0_write_write_3_stage_68;
  reg [31:0] bright_bright_update_0_write_write_3_stage_69;
  reg [31:0] bright_bright_update_0_write_write_3_stage_70;
  reg [31:0] bright_bright_update_0_write_write_3_stage_71;
  reg [31:0] bright_bright_update_0_write_write_3_stage_72;
  reg [31:0] bright_bright_update_0_write_write_3_stage_73;
  reg [31:0] bright_bright_update_0_write_write_3_stage_74;
  reg [31:0] bright_bright_update_0_write_write_3_stage_75;
  reg [31:0] bright_bright_update_0_write_write_3_stage_76;
  reg [31:0] bright_bright_update_0_write_write_3_stage_77;
  reg [31:0] bright_bright_update_0_write_write_3_stage_78;
  reg [31:0] bright_bright_update_0_write_write_3_stage_79;
  reg [31:0] bright_bright_update_0_write_write_3_stage_80;
  reg [31:0] bright_bright_update_0_write_write_3_stage_81;
  reg [31:0] bright_bright_update_0_write_write_3_stage_82;
  reg [31:0] bright_bright_update_0_write_write_3_stage_83;
  reg [31:0] bright_bright_update_0_write_write_3_stage_84;
  reg [31:0] bright_bright_update_0_write_write_3_stage_85;
  reg [31:0] bright_bright_update_0_write_write_3_stage_86;
  reg [31:0] bright_bright_update_0_write_write_3_stage_87;
  reg [31:0] bright_bright_update_0_write_write_3_stage_88;
  reg [31:0] bright_bright_update_0_write_write_3_stage_89;
  reg [31:0] bright_bright_update_0_write_write_3_stage_90;
  reg [31:0] bright_bright_update_0_write_write_3_stage_91;
  reg [31:0] bright_bright_update_0_write_write_3_stage_92;
  reg [31:0] bright_bright_update_0_write_write_3_stage_93;
  reg [31:0] bright_bright_update_0_write_write_3_stage_94;
  reg [31:0] bright_bright_update_0_write_write_3_stage_95;
  reg [31:0] bright_bright_update_0_write_write_3_stage_96;
  reg [31:0] bright_bright_update_0_write_write_3_stage_97;
  reg [31:0] bright_bright_update_0_write_write_3_stage_98;
  reg [31:0] bright_bright_update_0_write_write_3_stage_99;
  reg [31:0] bright_bright_update_0_write_write_3_stage_100;
  reg [31:0] bright_bright_update_0_write_write_3_stage_101;
  reg [31:0] bright_bright_update_0_write_write_3_stage_102;
  reg [31:0] bright_bright_update_0_write_write_3_stage_103;
  reg [31:0] bright_bright_update_0_write_write_3_stage_104;
  reg [31:0] bright_bright_update_0_write_write_3_stage_105;
  reg [31:0] bright_bright_update_0_write_write_3_stage_106;
  reg [31:0] bright_bright_update_0_write_write_3_stage_107;
  reg [31:0] bright_bright_update_0_write_write_3_stage_108;
  reg [31:0] bright_bright_update_0_write_write_3_stage_109;
  reg [31:0] bright_bright_update_0_write_write_3_stage_110;
  reg [31:0] bright_bright_update_0_write_write_3_stage_111;
  reg [31:0] bright_bright_update_0_write_write_3_stage_112;
  reg [31:0] bright_bright_update_0_write_write_3_stage_113;
  reg [31:0] bright_bright_update_0_write_write_3_stage_114;
  reg [31:0] bright_bright_update_0_write_write_3_stage_115;
  reg [31:0] bright_bright_update_0_write_write_3_stage_116;
  reg [31:0] bright_bright_update_0_write_write_3_stage_117;
  reg [31:0] bright_bright_update_0_write_write_3_stage_118;
  reg [31:0] bright_bright_update_0_write_write_3_stage_119;
  reg [31:0] bright_bright_update_0_write_write_3_stage_120;
  reg [31:0] bright_bright_update_0_write_write_3_stage_121;
  reg [31:0] bright_bright_update_0_write_write_3_stage_122;
  reg [31:0] bright_bright_update_0_write_write_3_stage_123;
  reg [31:0] bright_bright_update_0_write_write_3_stage_124;
  reg [31:0] bright_bright_update_0_write_write_3_stage_125;
  reg [31:0] bright_bright_update_0_write_write_3_stage_126;
  reg [31:0] bright_bright_update_0_write_write_3_stage_127;
  reg [31:0] bright_bright_update_0_write_write_3_stage_128;
  reg [31:0] bright_bright_update_0_write_write_3_stage_129;
  reg [31:0] bright_bright_update_0_write_write_3_stage_130;
  reg [31:0] bright_bright_update_0_write_write_3_stage_131;
  reg [31:0] bright_bright_update_0_write_write_3_stage_132;
  reg [31:0] bright_bright_update_0_write_write_3_stage_133;
  reg [31:0] bright_bright_update_0_write_write_3_stage_134;
  reg [31:0] bright_bright_update_0_write_write_3_stage_135;
  reg [31:0] bright_bright_update_0_write_write_3_stage_136;
  reg [31:0] bright_bright_update_0_write_write_3_stage_137;
  reg [31:0] bright_bright_update_0_write_write_3_stage_138;
  reg [31:0] bright_bright_update_0_write_write_3_stage_139;
  reg [31:0] bright_bright_update_0_write_write_3_stage_140;
  reg [31:0] bright_bright_update_0_write_write_3_stage_141;
  reg [31:0] bright_bright_update_0_write_write_3_stage_142;
  reg [31:0] bright_bright_update_0_write_write_3_stage_143;
  reg [31:0] bright_bright_update_0_write_write_3_stage_144;
  reg [31:0] bright_bright_update_0_write_write_3_stage_145;
  reg [31:0] bright_bright_update_0_write_write_3_stage_146;
  reg [31:0] bright_bright_update_0_write_write_3_stage_147;
  reg [31:0] bright_bright_update_0_write_write_3_stage_148;
  reg [31:0] bright_bright_update_0_write_write_3_stage_149;
  reg [31:0] bright_bright_update_0_write_write_3_stage_150;
  reg [31:0] bright_bright_update_0_write_write_3_stage_151;
  reg [31:0] bright_bright_update_0_write_write_3_stage_152;
  reg [31:0] bright_bright_update_0_write_write_3_stage_153;
  reg [31:0] bright_bright_update_0_write_write_3_stage_154;
  reg [31:0] bright_bright_update_0_write_write_3_stage_155;
  reg [31:0] bright_bright_update_0_write_write_3_stage_156;
  reg [31:0] bright_bright_update_0_write_write_3_stage_157;
  reg [31:0] bright_bright_update_0_write_write_3_stage_158;
  reg [31:0] bright_bright_update_0_write_write_3_stage_159;
  reg [31:0] bright_bright_update_0_write_write_3_stage_160;
  reg [31:0] bright_bright_update_0_write_write_3_stage_161;
  reg [31:0] bright_bright_update_0_write_write_3_stage_162;
  reg [31:0] bright_bright_update_0_write_write_3_stage_163;
  reg [31:0] bright_bright_update_0_write_write_3_stage_164;
  reg [31:0] bright_bright_update_0_write_write_3_stage_165;
  reg [31:0] bright_bright_update_0_write_write_3_stage_166;
  reg [31:0] bright_bright_update_0_write_write_3_stage_167;
  reg [31:0] bright_bright_update_0_write_write_3_stage_168;
  reg [31:0] bright_bright_update_0_write_write_3_stage_169;
  reg [31:0] bright_bright_update_0_write_write_3_stage_170;
  reg [31:0] bright_bright_update_0_write_write_3_stage_171;
  reg [31:0] bright_bright_update_0_write_write_3_stage_172;
  reg [31:0] bright_bright_update_0_write_write_3_stage_173;
  reg [31:0] bright_bright_update_0_write_write_3_stage_174;
  reg [31:0] bright_bright_update_0_write_write_3_stage_175;
  reg [31:0] bright_bright_update_0_write_write_3_stage_176;
  reg [31:0] bright_bright_update_0_write_write_3_stage_177;
  reg [31:0] bright_bright_update_0_write_write_3_stage_178;
  reg [31:0] bright_bright_update_0_write_write_3_stage_179;
  reg [31:0] bright_bright_update_0_write_write_3_stage_180;
  reg [31:0] bright_bright_update_0_write_write_3_stage_181;
  reg [31:0] in_dark_update_0_read_read_6_stage_11;
  reg [31:0] in_dark_update_0_read_read_6_stage_12;
  reg [31:0] in_dark_update_0_read_read_6_stage_13;
  reg [31:0] in_dark_update_0_read_read_6_stage_14;
  reg [31:0] in_dark_update_0_read_read_6_stage_15;
  reg [31:0] in_dark_update_0_read_read_6_stage_16;
  reg [31:0] in_dark_update_0_read_read_6_stage_17;
  reg [31:0] in_dark_update_0_read_read_6_stage_18;
  reg [31:0] in_dark_update_0_read_read_6_stage_19;
  reg [31:0] in_dark_update_0_read_read_6_stage_20;
  reg [31:0] in_dark_update_0_read_read_6_stage_21;
  reg [31:0] in_dark_update_0_read_read_6_stage_22;
  reg [31:0] in_dark_update_0_read_read_6_stage_23;
  reg [31:0] in_dark_update_0_read_read_6_stage_24;
  reg [31:0] in_dark_update_0_read_read_6_stage_25;
  reg [31:0] in_dark_update_0_read_read_6_stage_26;
  reg [31:0] in_dark_update_0_read_read_6_stage_27;
  reg [31:0] in_dark_update_0_read_read_6_stage_28;
  reg [31:0] in_dark_update_0_read_read_6_stage_29;
  reg [31:0] in_dark_update_0_read_read_6_stage_30;
  reg [31:0] in_dark_update_0_read_read_6_stage_31;
  reg [31:0] in_dark_update_0_read_read_6_stage_32;
  reg [31:0] in_dark_update_0_read_read_6_stage_33;
  reg [31:0] in_dark_update_0_read_read_6_stage_34;
  reg [31:0] in_dark_update_0_read_read_6_stage_35;
  reg [31:0] in_dark_update_0_read_read_6_stage_36;
  reg [31:0] in_dark_update_0_read_read_6_stage_37;
  reg [31:0] in_dark_update_0_read_read_6_stage_38;
  reg [31:0] in_dark_update_0_read_read_6_stage_39;
  reg [31:0] in_dark_update_0_read_read_6_stage_40;
  reg [31:0] in_dark_update_0_read_read_6_stage_41;
  reg [31:0] in_dark_update_0_read_read_6_stage_42;
  reg [31:0] in_dark_update_0_read_read_6_stage_43;
  reg [31:0] in_dark_update_0_read_read_6_stage_44;
  reg [31:0] in_dark_update_0_read_read_6_stage_45;
  reg [31:0] in_dark_update_0_read_read_6_stage_46;
  reg [31:0] in_dark_update_0_read_read_6_stage_47;
  reg [31:0] in_dark_update_0_read_read_6_stage_48;
  reg [31:0] in_dark_update_0_read_read_6_stage_49;
  reg [31:0] in_dark_update_0_read_read_6_stage_50;
  reg [31:0] in_dark_update_0_read_read_6_stage_51;
  reg [31:0] in_dark_update_0_read_read_6_stage_52;
  reg [31:0] in_dark_update_0_read_read_6_stage_53;
  reg [31:0] in_dark_update_0_read_read_6_stage_54;
  reg [31:0] in_dark_update_0_read_read_6_stage_55;
  reg [31:0] in_dark_update_0_read_read_6_stage_56;
  reg [31:0] in_dark_update_0_read_read_6_stage_57;
  reg [31:0] in_dark_update_0_read_read_6_stage_58;
  reg [31:0] in_dark_update_0_read_read_6_stage_59;
  reg [31:0] in_dark_update_0_read_read_6_stage_60;
  reg [31:0] in_dark_update_0_read_read_6_stage_61;
  reg [31:0] in_dark_update_0_read_read_6_stage_62;
  reg [31:0] in_dark_update_0_read_read_6_stage_63;
  reg [31:0] in_dark_update_0_read_read_6_stage_64;
  reg [31:0] in_dark_update_0_read_read_6_stage_65;
  reg [31:0] in_dark_update_0_read_read_6_stage_66;
  reg [31:0] in_dark_update_0_read_read_6_stage_67;
  reg [31:0] in_dark_update_0_read_read_6_stage_68;
  reg [31:0] in_dark_update_0_read_read_6_stage_69;
  reg [31:0] in_dark_update_0_read_read_6_stage_70;
  reg [31:0] in_dark_update_0_read_read_6_stage_71;
  reg [31:0] in_dark_update_0_read_read_6_stage_72;
  reg [31:0] in_dark_update_0_read_read_6_stage_73;
  reg [31:0] in_dark_update_0_read_read_6_stage_74;
  reg [31:0] in_dark_update_0_read_read_6_stage_75;
  reg [31:0] in_dark_update_0_read_read_6_stage_76;
  reg [31:0] in_dark_update_0_read_read_6_stage_77;
  reg [31:0] in_dark_update_0_read_read_6_stage_78;
  reg [31:0] in_dark_update_0_read_read_6_stage_79;
  reg [31:0] in_dark_update_0_read_read_6_stage_80;
  reg [31:0] in_dark_update_0_read_read_6_stage_81;
  reg [31:0] in_dark_update_0_read_read_6_stage_82;
  reg [31:0] in_dark_update_0_read_read_6_stage_83;
  reg [31:0] in_dark_update_0_read_read_6_stage_84;
  reg [31:0] in_dark_update_0_read_read_6_stage_85;
  reg [31:0] in_dark_update_0_read_read_6_stage_86;
  reg [31:0] in_dark_update_0_read_read_6_stage_87;
  reg [31:0] in_dark_update_0_read_read_6_stage_88;
  reg [31:0] in_dark_update_0_read_read_6_stage_89;
  reg [31:0] in_dark_update_0_read_read_6_stage_90;
  reg [31:0] in_dark_update_0_read_read_6_stage_91;
  reg [31:0] in_dark_update_0_read_read_6_stage_92;
  reg [31:0] in_dark_update_0_read_read_6_stage_93;
  reg [31:0] in_dark_update_0_read_read_6_stage_94;
  reg [31:0] in_dark_update_0_read_read_6_stage_95;
  reg [31:0] in_dark_update_0_read_read_6_stage_96;
  reg [31:0] in_dark_update_0_read_read_6_stage_97;
  reg [31:0] in_dark_update_0_read_read_6_stage_98;
  reg [31:0] in_dark_update_0_read_read_6_stage_99;
  reg [31:0] in_dark_update_0_read_read_6_stage_100;
  reg [31:0] in_dark_update_0_read_read_6_stage_101;
  reg [31:0] in_dark_update_0_read_read_6_stage_102;
  reg [31:0] in_dark_update_0_read_read_6_stage_103;
  reg [31:0] in_dark_update_0_read_read_6_stage_104;
  reg [31:0] in_dark_update_0_read_read_6_stage_105;
  reg [31:0] in_dark_update_0_read_read_6_stage_106;
  reg [31:0] in_dark_update_0_read_read_6_stage_107;
  reg [31:0] in_dark_update_0_read_read_6_stage_108;
  reg [31:0] in_dark_update_0_read_read_6_stage_109;
  reg [31:0] in_dark_update_0_read_read_6_stage_110;
  reg [31:0] in_dark_update_0_read_read_6_stage_111;
  reg [31:0] in_dark_update_0_read_read_6_stage_112;
  reg [31:0] in_dark_update_0_read_read_6_stage_113;
  reg [31:0] in_dark_update_0_read_read_6_stage_114;
  reg [31:0] in_dark_update_0_read_read_6_stage_115;
  reg [31:0] in_dark_update_0_read_read_6_stage_116;
  reg [31:0] in_dark_update_0_read_read_6_stage_117;
  reg [31:0] in_dark_update_0_read_read_6_stage_118;
  reg [31:0] in_dark_update_0_read_read_6_stage_119;
  reg [31:0] in_dark_update_0_read_read_6_stage_120;
  reg [31:0] in_dark_update_0_read_read_6_stage_121;
  reg [31:0] in_dark_update_0_read_read_6_stage_122;
  reg [31:0] in_dark_update_0_read_read_6_stage_123;
  reg [31:0] in_dark_update_0_read_read_6_stage_124;
  reg [31:0] in_dark_update_0_read_read_6_stage_125;
  reg [31:0] in_dark_update_0_read_read_6_stage_126;
  reg [31:0] in_dark_update_0_read_read_6_stage_127;
  reg [31:0] in_dark_update_0_read_read_6_stage_128;
  reg [31:0] in_dark_update_0_read_read_6_stage_129;
  reg [31:0] in_dark_update_0_read_read_6_stage_130;
  reg [31:0] in_dark_update_0_read_read_6_stage_131;
  reg [31:0] in_dark_update_0_read_read_6_stage_132;
  reg [31:0] in_dark_update_0_read_read_6_stage_133;
  reg [31:0] in_dark_update_0_read_read_6_stage_134;
  reg [31:0] in_dark_update_0_read_read_6_stage_135;
  reg [31:0] in_dark_update_0_read_read_6_stage_136;
  reg [31:0] in_dark_update_0_read_read_6_stage_137;
  reg [31:0] in_dark_update_0_read_read_6_stage_138;
  reg [31:0] in_dark_update_0_read_read_6_stage_139;
  reg [31:0] in_dark_update_0_read_read_6_stage_140;
  reg [31:0] in_dark_update_0_read_read_6_stage_141;
  reg [31:0] in_dark_update_0_read_read_6_stage_142;
  reg [31:0] in_dark_update_0_read_read_6_stage_143;
  reg [31:0] in_dark_update_0_read_read_6_stage_144;
  reg [31:0] in_dark_update_0_read_read_6_stage_145;
  reg [31:0] in_dark_update_0_read_read_6_stage_146;
  reg [31:0] in_dark_update_0_read_read_6_stage_147;
  reg [31:0] in_dark_update_0_read_read_6_stage_148;
  reg [31:0] in_dark_update_0_read_read_6_stage_149;
  reg [31:0] in_dark_update_0_read_read_6_stage_150;
  reg [31:0] in_dark_update_0_read_read_6_stage_151;
  reg [31:0] in_dark_update_0_read_read_6_stage_152;
  reg [31:0] in_dark_update_0_read_read_6_stage_153;
  reg [31:0] in_dark_update_0_read_read_6_stage_154;
  reg [31:0] in_dark_update_0_read_read_6_stage_155;
  reg [31:0] in_dark_update_0_read_read_6_stage_156;
  reg [31:0] in_dark_update_0_read_read_6_stage_157;
  reg [31:0] in_dark_update_0_read_read_6_stage_158;
  reg [31:0] in_dark_update_0_read_read_6_stage_159;
  reg [31:0] in_dark_update_0_read_read_6_stage_160;
  reg [31:0] in_dark_update_0_read_read_6_stage_161;
  reg [31:0] in_dark_update_0_read_read_6_stage_162;
  reg [31:0] in_dark_update_0_read_read_6_stage_163;
  reg [31:0] in_dark_update_0_read_read_6_stage_164;
  reg [31:0] in_dark_update_0_read_read_6_stage_165;
  reg [31:0] in_dark_update_0_read_read_6_stage_166;
  reg [31:0] in_dark_update_0_read_read_6_stage_167;
  reg [31:0] in_dark_update_0_read_read_6_stage_168;
  reg [31:0] in_dark_update_0_read_read_6_stage_169;
  reg [31:0] in_dark_update_0_read_read_6_stage_170;
  reg [31:0] in_dark_update_0_read_read_6_stage_171;
  reg [31:0] in_dark_update_0_read_read_6_stage_172;
  reg [31:0] in_dark_update_0_read_read_6_stage_173;
  reg [31:0] in_dark_update_0_read_read_6_stage_174;
  reg [31:0] in_dark_update_0_read_read_6_stage_175;
  reg [31:0] in_dark_update_0_read_read_6_stage_176;
  reg [31:0] in_dark_update_0_read_read_6_stage_177;
  reg [31:0] in_dark_update_0_read_read_6_stage_178;
  reg [31:0] in_dark_update_0_read_read_6_stage_179;
  reg [31:0] in_dark_update_0_read_read_6_stage_180;
  reg [31:0] in_dark_update_0_read_read_6_stage_181;
  reg [31:0] dark_update_0_stage_12;
  reg [31:0] dark_update_0_stage_13;
  reg [31:0] dark_update_0_stage_14;
  reg [31:0] dark_update_0_stage_15;
  reg [31:0] dark_update_0_stage_16;
  reg [31:0] dark_update_0_stage_17;
  reg [31:0] dark_update_0_stage_18;
  reg [31:0] dark_update_0_stage_19;
  reg [31:0] dark_update_0_stage_20;
  reg [31:0] dark_update_0_stage_21;
  reg [31:0] dark_update_0_stage_22;
  reg [31:0] dark_update_0_stage_23;
  reg [31:0] dark_update_0_stage_24;
  reg [31:0] dark_update_0_stage_25;
  reg [31:0] dark_update_0_stage_26;
  reg [31:0] dark_update_0_stage_27;
  reg [31:0] dark_update_0_stage_28;
  reg [31:0] dark_update_0_stage_29;
  reg [31:0] dark_update_0_stage_30;
  reg [31:0] dark_update_0_stage_31;
  reg [31:0] dark_update_0_stage_32;
  reg [31:0] dark_update_0_stage_33;
  reg [31:0] dark_update_0_stage_34;
  reg [31:0] dark_update_0_stage_35;
  reg [31:0] dark_update_0_stage_36;
  reg [31:0] dark_update_0_stage_37;
  reg [31:0] dark_update_0_stage_38;
  reg [31:0] dark_update_0_stage_39;
  reg [31:0] dark_update_0_stage_40;
  reg [31:0] dark_update_0_stage_41;
  reg [31:0] dark_update_0_stage_42;
  reg [31:0] dark_update_0_stage_43;
  reg [31:0] dark_update_0_stage_44;
  reg [31:0] dark_update_0_stage_45;
  reg [31:0] dark_update_0_stage_46;
  reg [31:0] dark_update_0_stage_47;
  reg [31:0] dark_update_0_stage_48;
  reg [31:0] dark_update_0_stage_49;
  reg [31:0] dark_update_0_stage_50;
  reg [31:0] dark_update_0_stage_51;
  reg [31:0] dark_update_0_stage_52;
  reg [31:0] dark_update_0_stage_53;
  reg [31:0] dark_update_0_stage_54;
  reg [31:0] dark_update_0_stage_55;
  reg [31:0] dark_update_0_stage_56;
  reg [31:0] dark_update_0_stage_57;
  reg [31:0] dark_update_0_stage_58;
  reg [31:0] dark_update_0_stage_59;
  reg [31:0] dark_update_0_stage_60;
  reg [31:0] dark_update_0_stage_61;
  reg [31:0] dark_update_0_stage_62;
  reg [31:0] dark_update_0_stage_63;
  reg [31:0] dark_update_0_stage_64;
  reg [31:0] dark_update_0_stage_65;
  reg [31:0] dark_update_0_stage_66;
  reg [31:0] dark_update_0_stage_67;
  reg [31:0] dark_update_0_stage_68;
  reg [31:0] dark_update_0_stage_69;
  reg [31:0] dark_update_0_stage_70;
  reg [31:0] dark_update_0_stage_71;
  reg [31:0] dark_update_0_stage_72;
  reg [31:0] dark_update_0_stage_73;
  reg [31:0] dark_update_0_stage_74;
  reg [31:0] dark_update_0_stage_75;
  reg [31:0] dark_update_0_stage_76;
  reg [31:0] dark_update_0_stage_77;
  reg [31:0] dark_update_0_stage_78;
  reg [31:0] dark_update_0_stage_79;
  reg [31:0] dark_update_0_stage_80;
  reg [31:0] dark_update_0_stage_81;
  reg [31:0] dark_update_0_stage_82;
  reg [31:0] dark_update_0_stage_83;
  reg [31:0] dark_update_0_stage_84;
  reg [31:0] dark_update_0_stage_85;
  reg [31:0] dark_update_0_stage_86;
  reg [31:0] dark_update_0_stage_87;
  reg [31:0] dark_update_0_stage_88;
  reg [31:0] dark_update_0_stage_89;
  reg [31:0] dark_update_0_stage_90;
  reg [31:0] dark_update_0_stage_91;
  reg [31:0] dark_update_0_stage_92;
  reg [31:0] dark_update_0_stage_93;
  reg [31:0] dark_update_0_stage_94;
  reg [31:0] dark_update_0_stage_95;
  reg [31:0] dark_update_0_stage_96;
  reg [31:0] dark_update_0_stage_97;
  reg [31:0] dark_update_0_stage_98;
  reg [31:0] dark_update_0_stage_99;
  reg [31:0] dark_update_0_stage_100;
  reg [31:0] dark_update_0_stage_101;
  reg [31:0] dark_update_0_stage_102;
  reg [31:0] dark_update_0_stage_103;
  reg [31:0] dark_update_0_stage_104;
  reg [31:0] dark_update_0_stage_105;
  reg [31:0] dark_update_0_stage_106;
  reg [31:0] dark_update_0_stage_107;
  reg [31:0] dark_update_0_stage_108;
  reg [31:0] dark_update_0_stage_109;
  reg [31:0] dark_update_0_stage_110;
  reg [31:0] dark_update_0_stage_111;
  reg [31:0] dark_update_0_stage_112;
  reg [31:0] dark_update_0_stage_113;
  reg [31:0] dark_update_0_stage_114;
  reg [31:0] dark_update_0_stage_115;
  reg [31:0] dark_update_0_stage_116;
  reg [31:0] dark_update_0_stage_117;
  reg [31:0] dark_update_0_stage_118;
  reg [31:0] dark_update_0_stage_119;
  reg [31:0] dark_update_0_stage_120;
  reg [31:0] dark_update_0_stage_121;
  reg [31:0] dark_update_0_stage_122;
  reg [31:0] dark_update_0_stage_123;
  reg [31:0] dark_update_0_stage_124;
  reg [31:0] dark_update_0_stage_125;
  reg [31:0] dark_update_0_stage_126;
  reg [31:0] dark_update_0_stage_127;
  reg [31:0] dark_update_0_stage_128;
  reg [31:0] dark_update_0_stage_129;
  reg [31:0] dark_update_0_stage_130;
  reg [31:0] dark_update_0_stage_131;
  reg [31:0] dark_update_0_stage_132;
  reg [31:0] dark_update_0_stage_133;
  reg [31:0] dark_update_0_stage_134;
  reg [31:0] dark_update_0_stage_135;
  reg [31:0] dark_update_0_stage_136;
  reg [31:0] dark_update_0_stage_137;
  reg [31:0] dark_update_0_stage_138;
  reg [31:0] dark_update_0_stage_139;
  reg [31:0] dark_update_0_stage_140;
  reg [31:0] dark_update_0_stage_141;
  reg [31:0] dark_update_0_stage_142;
  reg [31:0] dark_update_0_stage_143;
  reg [31:0] dark_update_0_stage_144;
  reg [31:0] dark_update_0_stage_145;
  reg [31:0] dark_update_0_stage_146;
  reg [31:0] dark_update_0_stage_147;
  reg [31:0] dark_update_0_stage_148;
  reg [31:0] dark_update_0_stage_149;
  reg [31:0] dark_update_0_stage_150;
  reg [31:0] dark_update_0_stage_151;
  reg [31:0] dark_update_0_stage_152;
  reg [31:0] dark_update_0_stage_153;
  reg [31:0] dark_update_0_stage_154;
  reg [31:0] dark_update_0_stage_155;
  reg [31:0] dark_update_0_stage_156;
  reg [31:0] dark_update_0_stage_157;
  reg [31:0] dark_update_0_stage_158;
  reg [31:0] dark_update_0_stage_159;
  reg [31:0] dark_update_0_stage_160;
  reg [31:0] dark_update_0_stage_161;
  reg [31:0] dark_update_0_stage_162;
  reg [31:0] dark_update_0_stage_163;
  reg [31:0] dark_update_0_stage_164;
  reg [31:0] dark_update_0_stage_165;
  reg [31:0] dark_update_0_stage_166;
  reg [31:0] dark_update_0_stage_167;
  reg [31:0] dark_update_0_stage_168;
  reg [31:0] dark_update_0_stage_169;
  reg [31:0] dark_update_0_stage_170;
  reg [31:0] dark_update_0_stage_171;
  reg [31:0] dark_update_0_stage_172;
  reg [31:0] dark_update_0_stage_173;
  reg [31:0] dark_update_0_stage_174;
  reg [31:0] dark_update_0_stage_175;
  reg [31:0] dark_update_0_stage_176;
  reg [31:0] dark_update_0_stage_177;
  reg [31:0] dark_update_0_stage_178;
  reg [31:0] dark_update_0_stage_179;
  reg [31:0] dark_update_0_stage_180;
  reg [31:0] dark_update_0_stage_181;
  reg [31:0] dark_dark_update_0_write_write_7_stage_13;
  reg [31:0] dark_dark_update_0_write_write_7_stage_14;
  reg [31:0] dark_dark_update_0_write_write_7_stage_15;
  reg [31:0] dark_dark_update_0_write_write_7_stage_16;
  reg [31:0] dark_dark_update_0_write_write_7_stage_17;
  reg [31:0] dark_dark_update_0_write_write_7_stage_18;
  reg [31:0] dark_dark_update_0_write_write_7_stage_19;
  reg [31:0] dark_dark_update_0_write_write_7_stage_20;
  reg [31:0] dark_dark_update_0_write_write_7_stage_21;
  reg [31:0] dark_dark_update_0_write_write_7_stage_22;
  reg [31:0] dark_dark_update_0_write_write_7_stage_23;
  reg [31:0] dark_dark_update_0_write_write_7_stage_24;
  reg [31:0] dark_dark_update_0_write_write_7_stage_25;
  reg [31:0] dark_dark_update_0_write_write_7_stage_26;
  reg [31:0] dark_dark_update_0_write_write_7_stage_27;
  reg [31:0] dark_dark_update_0_write_write_7_stage_28;
  reg [31:0] dark_dark_update_0_write_write_7_stage_29;
  reg [31:0] dark_dark_update_0_write_write_7_stage_30;
  reg [31:0] dark_dark_update_0_write_write_7_stage_31;
  reg [31:0] dark_dark_update_0_write_write_7_stage_32;
  reg [31:0] dark_dark_update_0_write_write_7_stage_33;
  reg [31:0] dark_dark_update_0_write_write_7_stage_34;
  reg [31:0] dark_dark_update_0_write_write_7_stage_35;
  reg [31:0] dark_dark_update_0_write_write_7_stage_36;
  reg [31:0] dark_dark_update_0_write_write_7_stage_37;
  reg [31:0] dark_dark_update_0_write_write_7_stage_38;
  reg [31:0] dark_dark_update_0_write_write_7_stage_39;
  reg [31:0] dark_dark_update_0_write_write_7_stage_40;
  reg [31:0] dark_dark_update_0_write_write_7_stage_41;
  reg [31:0] dark_dark_update_0_write_write_7_stage_42;
  reg [31:0] dark_dark_update_0_write_write_7_stage_43;
  reg [31:0] dark_dark_update_0_write_write_7_stage_44;
  reg [31:0] dark_dark_update_0_write_write_7_stage_45;
  reg [31:0] dark_dark_update_0_write_write_7_stage_46;
  reg [31:0] dark_dark_update_0_write_write_7_stage_47;
  reg [31:0] dark_dark_update_0_write_write_7_stage_48;
  reg [31:0] dark_dark_update_0_write_write_7_stage_49;
  reg [31:0] dark_dark_update_0_write_write_7_stage_50;
  reg [31:0] dark_dark_update_0_write_write_7_stage_51;
  reg [31:0] dark_dark_update_0_write_write_7_stage_52;
  reg [31:0] dark_dark_update_0_write_write_7_stage_53;
  reg [31:0] dark_dark_update_0_write_write_7_stage_54;
  reg [31:0] dark_dark_update_0_write_write_7_stage_55;
  reg [31:0] dark_dark_update_0_write_write_7_stage_56;
  reg [31:0] dark_dark_update_0_write_write_7_stage_57;
  reg [31:0] dark_dark_update_0_write_write_7_stage_58;
  reg [31:0] dark_dark_update_0_write_write_7_stage_59;
  reg [31:0] dark_dark_update_0_write_write_7_stage_60;
  reg [31:0] dark_dark_update_0_write_write_7_stage_61;
  reg [31:0] dark_dark_update_0_write_write_7_stage_62;
  reg [31:0] dark_dark_update_0_write_write_7_stage_63;
  reg [31:0] dark_dark_update_0_write_write_7_stage_64;
  reg [31:0] dark_dark_update_0_write_write_7_stage_65;
  reg [31:0] dark_dark_update_0_write_write_7_stage_66;
  reg [31:0] dark_dark_update_0_write_write_7_stage_67;
  reg [31:0] dark_dark_update_0_write_write_7_stage_68;
  reg [31:0] dark_dark_update_0_write_write_7_stage_69;
  reg [31:0] dark_dark_update_0_write_write_7_stage_70;
  reg [31:0] dark_dark_update_0_write_write_7_stage_71;
  reg [31:0] dark_dark_update_0_write_write_7_stage_72;
  reg [31:0] dark_dark_update_0_write_write_7_stage_73;
  reg [31:0] dark_dark_update_0_write_write_7_stage_74;
  reg [31:0] dark_dark_update_0_write_write_7_stage_75;
  reg [31:0] dark_dark_update_0_write_write_7_stage_76;
  reg [31:0] dark_dark_update_0_write_write_7_stage_77;
  reg [31:0] dark_dark_update_0_write_write_7_stage_78;
  reg [31:0] dark_dark_update_0_write_write_7_stage_79;
  reg [31:0] dark_dark_update_0_write_write_7_stage_80;
  reg [31:0] dark_dark_update_0_write_write_7_stage_81;
  reg [31:0] dark_dark_update_0_write_write_7_stage_82;
  reg [31:0] dark_dark_update_0_write_write_7_stage_83;
  reg [31:0] dark_dark_update_0_write_write_7_stage_84;
  reg [31:0] dark_dark_update_0_write_write_7_stage_85;
  reg [31:0] dark_dark_update_0_write_write_7_stage_86;
  reg [31:0] dark_dark_update_0_write_write_7_stage_87;
  reg [31:0] dark_dark_update_0_write_write_7_stage_88;
  reg [31:0] dark_dark_update_0_write_write_7_stage_89;
  reg [31:0] dark_dark_update_0_write_write_7_stage_90;
  reg [31:0] dark_dark_update_0_write_write_7_stage_91;
  reg [31:0] dark_dark_update_0_write_write_7_stage_92;
  reg [31:0] dark_dark_update_0_write_write_7_stage_93;
  reg [31:0] dark_dark_update_0_write_write_7_stage_94;
  reg [31:0] dark_dark_update_0_write_write_7_stage_95;
  reg [31:0] dark_dark_update_0_write_write_7_stage_96;
  reg [31:0] dark_dark_update_0_write_write_7_stage_97;
  reg [31:0] dark_dark_update_0_write_write_7_stage_98;
  reg [31:0] dark_dark_update_0_write_write_7_stage_99;
  reg [31:0] dark_dark_update_0_write_write_7_stage_100;
  reg [31:0] dark_dark_update_0_write_write_7_stage_101;
  reg [31:0] dark_dark_update_0_write_write_7_stage_102;
  reg [31:0] dark_dark_update_0_write_write_7_stage_103;
  reg [31:0] dark_dark_update_0_write_write_7_stage_104;
  reg [31:0] dark_dark_update_0_write_write_7_stage_105;
  reg [31:0] dark_dark_update_0_write_write_7_stage_106;
  reg [31:0] dark_dark_update_0_write_write_7_stage_107;
  reg [31:0] dark_dark_update_0_write_write_7_stage_108;
  reg [31:0] dark_dark_update_0_write_write_7_stage_109;
  reg [31:0] dark_dark_update_0_write_write_7_stage_110;
  reg [31:0] dark_dark_update_0_write_write_7_stage_111;
  reg [31:0] dark_dark_update_0_write_write_7_stage_112;
  reg [31:0] dark_dark_update_0_write_write_7_stage_113;
  reg [31:0] dark_dark_update_0_write_write_7_stage_114;
  reg [31:0] dark_dark_update_0_write_write_7_stage_115;
  reg [31:0] dark_dark_update_0_write_write_7_stage_116;
  reg [31:0] dark_dark_update_0_write_write_7_stage_117;
  reg [31:0] dark_dark_update_0_write_write_7_stage_118;
  reg [31:0] dark_dark_update_0_write_write_7_stage_119;
  reg [31:0] dark_dark_update_0_write_write_7_stage_120;
  reg [31:0] dark_dark_update_0_write_write_7_stage_121;
  reg [31:0] dark_dark_update_0_write_write_7_stage_122;
  reg [31:0] dark_dark_update_0_write_write_7_stage_123;
  reg [31:0] dark_dark_update_0_write_write_7_stage_124;
  reg [31:0] dark_dark_update_0_write_write_7_stage_125;
  reg [31:0] dark_dark_update_0_write_write_7_stage_126;
  reg [31:0] dark_dark_update_0_write_write_7_stage_127;
  reg [31:0] dark_dark_update_0_write_write_7_stage_128;
  reg [31:0] dark_dark_update_0_write_write_7_stage_129;
  reg [31:0] dark_dark_update_0_write_write_7_stage_130;
  reg [31:0] dark_dark_update_0_write_write_7_stage_131;
  reg [31:0] dark_dark_update_0_write_write_7_stage_132;
  reg [31:0] dark_dark_update_0_write_write_7_stage_133;
  reg [31:0] dark_dark_update_0_write_write_7_stage_134;
  reg [31:0] dark_dark_update_0_write_write_7_stage_135;
  reg [31:0] dark_dark_update_0_write_write_7_stage_136;
  reg [31:0] dark_dark_update_0_write_write_7_stage_137;
  reg [31:0] dark_dark_update_0_write_write_7_stage_138;
  reg [31:0] dark_dark_update_0_write_write_7_stage_139;
  reg [31:0] dark_dark_update_0_write_write_7_stage_140;
  reg [31:0] dark_dark_update_0_write_write_7_stage_141;
  reg [31:0] dark_dark_update_0_write_write_7_stage_142;
  reg [31:0] dark_dark_update_0_write_write_7_stage_143;
  reg [31:0] dark_dark_update_0_write_write_7_stage_144;
  reg [31:0] dark_dark_update_0_write_write_7_stage_145;
  reg [31:0] dark_dark_update_0_write_write_7_stage_146;
  reg [31:0] dark_dark_update_0_write_write_7_stage_147;
  reg [31:0] dark_dark_update_0_write_write_7_stage_148;
  reg [31:0] dark_dark_update_0_write_write_7_stage_149;
  reg [31:0] dark_dark_update_0_write_write_7_stage_150;
  reg [31:0] dark_dark_update_0_write_write_7_stage_151;
  reg [31:0] dark_dark_update_0_write_write_7_stage_152;
  reg [31:0] dark_dark_update_0_write_write_7_stage_153;
  reg [31:0] dark_dark_update_0_write_write_7_stage_154;
  reg [31:0] dark_dark_update_0_write_write_7_stage_155;
  reg [31:0] dark_dark_update_0_write_write_7_stage_156;
  reg [31:0] dark_dark_update_0_write_write_7_stage_157;
  reg [31:0] dark_dark_update_0_write_write_7_stage_158;
  reg [31:0] dark_dark_update_0_write_write_7_stage_159;
  reg [31:0] dark_dark_update_0_write_write_7_stage_160;
  reg [31:0] dark_dark_update_0_write_write_7_stage_161;
  reg [31:0] dark_dark_update_0_write_write_7_stage_162;
  reg [31:0] dark_dark_update_0_write_write_7_stage_163;
  reg [31:0] dark_dark_update_0_write_write_7_stage_164;
  reg [31:0] dark_dark_update_0_write_write_7_stage_165;
  reg [31:0] dark_dark_update_0_write_write_7_stage_166;
  reg [31:0] dark_dark_update_0_write_write_7_stage_167;
  reg [31:0] dark_dark_update_0_write_write_7_stage_168;
  reg [31:0] dark_dark_update_0_write_write_7_stage_169;
  reg [31:0] dark_dark_update_0_write_write_7_stage_170;
  reg [31:0] dark_dark_update_0_write_write_7_stage_171;
  reg [31:0] dark_dark_update_0_write_write_7_stage_172;
  reg [31:0] dark_dark_update_0_write_write_7_stage_173;
  reg [31:0] dark_dark_update_0_write_write_7_stage_174;
  reg [31:0] dark_dark_update_0_write_write_7_stage_175;
  reg [31:0] dark_dark_update_0_write_write_7_stage_176;
  reg [31:0] dark_dark_update_0_write_write_7_stage_177;
  reg [31:0] dark_dark_update_0_write_write_7_stage_178;
  reg [31:0] dark_dark_update_0_write_write_7_stage_179;
  reg [31:0] dark_dark_update_0_write_write_7_stage_180;
  reg [31:0] dark_dark_update_0_write_write_7_stage_181;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_17;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_18;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_19;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_20;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_21;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_22;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_23;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_24;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_25;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_26;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_27;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_28;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_29;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_30;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_31;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_32;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_33;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_34;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_35;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_36;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_37;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_38;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_39;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_40;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_41;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_42;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_43;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_44;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_45;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_46;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_47;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_48;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_49;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_50;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_51;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_52;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_53;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_54;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_55;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_56;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_57;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_58;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_59;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_60;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_61;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_62;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_63;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_64;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_65;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_66;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_67;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_68;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_69;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_70;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_71;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_72;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_73;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_74;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_75;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_76;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_77;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_78;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_79;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_80;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_81;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_82;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_83;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_84;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_85;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_86;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_87;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_88;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_89;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_90;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_91;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_92;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_93;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_94;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_95;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_96;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_97;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_98;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_99;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_100;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_101;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_102;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_103;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_104;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_105;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_106;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_107;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_108;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_109;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_110;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_111;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_112;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_113;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_114;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_115;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_116;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_117;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_118;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_119;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_120;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_121;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_122;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_123;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_124;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_125;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_126;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_127;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_128;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_129;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_130;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_131;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_132;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_133;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_134;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_135;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_136;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_137;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_138;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_139;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_140;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_141;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_142;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_143;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_144;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_145;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_146;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_147;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_148;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_149;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_150;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_151;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_152;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_153;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_154;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_155;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_156;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_157;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_158;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_159;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_160;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_161;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_162;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_163;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_164;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_165;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_166;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_167;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_168;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_169;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_170;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_171;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_172;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_173;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_174;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_175;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_176;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_177;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_178;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_179;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_180;
  reg [287:0] dark_dark_gauss_blur_1_update_0_read_read_10_stage_181;
  reg [31:0] dark_gauss_blur_1_update_0_stage_18;
  reg [31:0] dark_gauss_blur_1_update_0_stage_19;
  reg [31:0] dark_gauss_blur_1_update_0_stage_20;
  reg [31:0] dark_gauss_blur_1_update_0_stage_21;
  reg [31:0] dark_gauss_blur_1_update_0_stage_22;
  reg [31:0] dark_gauss_blur_1_update_0_stage_23;
  reg [31:0] dark_gauss_blur_1_update_0_stage_24;
  reg [31:0] dark_gauss_blur_1_update_0_stage_25;
  reg [31:0] dark_gauss_blur_1_update_0_stage_26;
  reg [31:0] dark_gauss_blur_1_update_0_stage_27;
  reg [31:0] dark_gauss_blur_1_update_0_stage_28;
  reg [31:0] dark_gauss_blur_1_update_0_stage_29;
  reg [31:0] dark_gauss_blur_1_update_0_stage_30;
  reg [31:0] dark_gauss_blur_1_update_0_stage_31;
  reg [31:0] dark_gauss_blur_1_update_0_stage_32;
  reg [31:0] dark_gauss_blur_1_update_0_stage_33;
  reg [31:0] dark_gauss_blur_1_update_0_stage_34;
  reg [31:0] dark_gauss_blur_1_update_0_stage_35;
  reg [31:0] dark_gauss_blur_1_update_0_stage_36;
  reg [31:0] dark_gauss_blur_1_update_0_stage_37;
  reg [31:0] dark_gauss_blur_1_update_0_stage_38;
  reg [31:0] dark_gauss_blur_1_update_0_stage_39;
  reg [31:0] dark_gauss_blur_1_update_0_stage_40;
  reg [31:0] dark_gauss_blur_1_update_0_stage_41;
  reg [31:0] dark_gauss_blur_1_update_0_stage_42;
  reg [31:0] dark_gauss_blur_1_update_0_stage_43;
  reg [31:0] dark_gauss_blur_1_update_0_stage_44;
  reg [31:0] dark_gauss_blur_1_update_0_stage_45;
  reg [31:0] dark_gauss_blur_1_update_0_stage_46;
  reg [31:0] dark_gauss_blur_1_update_0_stage_47;
  reg [31:0] dark_gauss_blur_1_update_0_stage_48;
  reg [31:0] dark_gauss_blur_1_update_0_stage_49;
  reg [31:0] dark_gauss_blur_1_update_0_stage_50;
  reg [31:0] dark_gauss_blur_1_update_0_stage_51;
  reg [31:0] dark_gauss_blur_1_update_0_stage_52;
  reg [31:0] dark_gauss_blur_1_update_0_stage_53;
  reg [31:0] dark_gauss_blur_1_update_0_stage_54;
  reg [31:0] dark_gauss_blur_1_update_0_stage_55;
  reg [31:0] dark_gauss_blur_1_update_0_stage_56;
  reg [31:0] dark_gauss_blur_1_update_0_stage_57;
  reg [31:0] dark_gauss_blur_1_update_0_stage_58;
  reg [31:0] dark_gauss_blur_1_update_0_stage_59;
  reg [31:0] dark_gauss_blur_1_update_0_stage_60;
  reg [31:0] dark_gauss_blur_1_update_0_stage_61;
  reg [31:0] dark_gauss_blur_1_update_0_stage_62;
  reg [31:0] dark_gauss_blur_1_update_0_stage_63;
  reg [31:0] dark_gauss_blur_1_update_0_stage_64;
  reg [31:0] dark_gauss_blur_1_update_0_stage_65;
  reg [31:0] dark_gauss_blur_1_update_0_stage_66;
  reg [31:0] dark_gauss_blur_1_update_0_stage_67;
  reg [31:0] dark_gauss_blur_1_update_0_stage_68;
  reg [31:0] dark_gauss_blur_1_update_0_stage_69;
  reg [31:0] dark_gauss_blur_1_update_0_stage_70;
  reg [31:0] dark_gauss_blur_1_update_0_stage_71;
  reg [31:0] dark_gauss_blur_1_update_0_stage_72;
  reg [31:0] dark_gauss_blur_1_update_0_stage_73;
  reg [31:0] dark_gauss_blur_1_update_0_stage_74;
  reg [31:0] dark_gauss_blur_1_update_0_stage_75;
  reg [31:0] dark_gauss_blur_1_update_0_stage_76;
  reg [31:0] dark_gauss_blur_1_update_0_stage_77;
  reg [31:0] dark_gauss_blur_1_update_0_stage_78;
  reg [31:0] dark_gauss_blur_1_update_0_stage_79;
  reg [31:0] dark_gauss_blur_1_update_0_stage_80;
  reg [31:0] dark_gauss_blur_1_update_0_stage_81;
  reg [31:0] dark_gauss_blur_1_update_0_stage_82;
  reg [31:0] dark_gauss_blur_1_update_0_stage_83;
  reg [31:0] dark_gauss_blur_1_update_0_stage_84;
  reg [31:0] dark_gauss_blur_1_update_0_stage_85;
  reg [31:0] dark_gauss_blur_1_update_0_stage_86;
  reg [31:0] dark_gauss_blur_1_update_0_stage_87;
  reg [31:0] dark_gauss_blur_1_update_0_stage_88;
  reg [31:0] dark_gauss_blur_1_update_0_stage_89;
  reg [31:0] dark_gauss_blur_1_update_0_stage_90;
  reg [31:0] dark_gauss_blur_1_update_0_stage_91;
  reg [31:0] dark_gauss_blur_1_update_0_stage_92;
  reg [31:0] dark_gauss_blur_1_update_0_stage_93;
  reg [31:0] dark_gauss_blur_1_update_0_stage_94;
  reg [31:0] dark_gauss_blur_1_update_0_stage_95;
  reg [31:0] dark_gauss_blur_1_update_0_stage_96;
  reg [31:0] dark_gauss_blur_1_update_0_stage_97;
  reg [31:0] dark_gauss_blur_1_update_0_stage_98;
  reg [31:0] dark_gauss_blur_1_update_0_stage_99;
  reg [31:0] dark_gauss_blur_1_update_0_stage_100;
  reg [31:0] dark_gauss_blur_1_update_0_stage_101;
  reg [31:0] dark_gauss_blur_1_update_0_stage_102;
  reg [31:0] dark_gauss_blur_1_update_0_stage_103;
  reg [31:0] dark_gauss_blur_1_update_0_stage_104;
  reg [31:0] dark_gauss_blur_1_update_0_stage_105;
  reg [31:0] dark_gauss_blur_1_update_0_stage_106;
  reg [31:0] dark_gauss_blur_1_update_0_stage_107;
  reg [31:0] dark_gauss_blur_1_update_0_stage_108;
  reg [31:0] dark_gauss_blur_1_update_0_stage_109;
  reg [31:0] dark_gauss_blur_1_update_0_stage_110;
  reg [31:0] dark_gauss_blur_1_update_0_stage_111;
  reg [31:0] dark_gauss_blur_1_update_0_stage_112;
  reg [31:0] dark_gauss_blur_1_update_0_stage_113;
  reg [31:0] dark_gauss_blur_1_update_0_stage_114;
  reg [31:0] dark_gauss_blur_1_update_0_stage_115;
  reg [31:0] dark_gauss_blur_1_update_0_stage_116;
  reg [31:0] dark_gauss_blur_1_update_0_stage_117;
  reg [31:0] dark_gauss_blur_1_update_0_stage_118;
  reg [31:0] dark_gauss_blur_1_update_0_stage_119;
  reg [31:0] dark_gauss_blur_1_update_0_stage_120;
  reg [31:0] dark_gauss_blur_1_update_0_stage_121;
  reg [31:0] dark_gauss_blur_1_update_0_stage_122;
  reg [31:0] dark_gauss_blur_1_update_0_stage_123;
  reg [31:0] dark_gauss_blur_1_update_0_stage_124;
  reg [31:0] dark_gauss_blur_1_update_0_stage_125;
  reg [31:0] dark_gauss_blur_1_update_0_stage_126;
  reg [31:0] dark_gauss_blur_1_update_0_stage_127;
  reg [31:0] dark_gauss_blur_1_update_0_stage_128;
  reg [31:0] dark_gauss_blur_1_update_0_stage_129;
  reg [31:0] dark_gauss_blur_1_update_0_stage_130;
  reg [31:0] dark_gauss_blur_1_update_0_stage_131;
  reg [31:0] dark_gauss_blur_1_update_0_stage_132;
  reg [31:0] dark_gauss_blur_1_update_0_stage_133;
  reg [31:0] dark_gauss_blur_1_update_0_stage_134;
  reg [31:0] dark_gauss_blur_1_update_0_stage_135;
  reg [31:0] dark_gauss_blur_1_update_0_stage_136;
  reg [31:0] dark_gauss_blur_1_update_0_stage_137;
  reg [31:0] dark_gauss_blur_1_update_0_stage_138;
  reg [31:0] dark_gauss_blur_1_update_0_stage_139;
  reg [31:0] dark_gauss_blur_1_update_0_stage_140;
  reg [31:0] dark_gauss_blur_1_update_0_stage_141;
  reg [31:0] dark_gauss_blur_1_update_0_stage_142;
  reg [31:0] dark_gauss_blur_1_update_0_stage_143;
  reg [31:0] dark_gauss_blur_1_update_0_stage_144;
  reg [31:0] dark_gauss_blur_1_update_0_stage_145;
  reg [31:0] dark_gauss_blur_1_update_0_stage_146;
  reg [31:0] dark_gauss_blur_1_update_0_stage_147;
  reg [31:0] dark_gauss_blur_1_update_0_stage_148;
  reg [31:0] dark_gauss_blur_1_update_0_stage_149;
  reg [31:0] dark_gauss_blur_1_update_0_stage_150;
  reg [31:0] dark_gauss_blur_1_update_0_stage_151;
  reg [31:0] dark_gauss_blur_1_update_0_stage_152;
  reg [31:0] dark_gauss_blur_1_update_0_stage_153;
  reg [31:0] dark_gauss_blur_1_update_0_stage_154;
  reg [31:0] dark_gauss_blur_1_update_0_stage_155;
  reg [31:0] dark_gauss_blur_1_update_0_stage_156;
  reg [31:0] dark_gauss_blur_1_update_0_stage_157;
  reg [31:0] dark_gauss_blur_1_update_0_stage_158;
  reg [31:0] dark_gauss_blur_1_update_0_stage_159;
  reg [31:0] dark_gauss_blur_1_update_0_stage_160;
  reg [31:0] dark_gauss_blur_1_update_0_stage_161;
  reg [31:0] dark_gauss_blur_1_update_0_stage_162;
  reg [31:0] dark_gauss_blur_1_update_0_stage_163;
  reg [31:0] dark_gauss_blur_1_update_0_stage_164;
  reg [31:0] dark_gauss_blur_1_update_0_stage_165;
  reg [31:0] dark_gauss_blur_1_update_0_stage_166;
  reg [31:0] dark_gauss_blur_1_update_0_stage_167;
  reg [31:0] dark_gauss_blur_1_update_0_stage_168;
  reg [31:0] dark_gauss_blur_1_update_0_stage_169;
  reg [31:0] dark_gauss_blur_1_update_0_stage_170;
  reg [31:0] dark_gauss_blur_1_update_0_stage_171;
  reg [31:0] dark_gauss_blur_1_update_0_stage_172;
  reg [31:0] dark_gauss_blur_1_update_0_stage_173;
  reg [31:0] dark_gauss_blur_1_update_0_stage_174;
  reg [31:0] dark_gauss_blur_1_update_0_stage_175;
  reg [31:0] dark_gauss_blur_1_update_0_stage_176;
  reg [31:0] dark_gauss_blur_1_update_0_stage_177;
  reg [31:0] dark_gauss_blur_1_update_0_stage_178;
  reg [31:0] dark_gauss_blur_1_update_0_stage_179;
  reg [31:0] dark_gauss_blur_1_update_0_stage_180;
  reg [31:0] dark_gauss_blur_1_update_0_stage_181;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_60;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_61;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_62;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_63;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_64;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_65;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_66;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_67;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_68;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_69;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_70;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_71;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_72;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_73;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_74;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_75;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_76;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_77;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_78;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_79;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_80;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_81;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_82;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_83;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_84;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_85;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_86;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_87;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_88;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_89;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_90;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_91;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_92;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_93;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_94;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_95;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_96;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_97;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_98;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_99;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_100;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_101;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_102;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_103;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_104;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_105;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_106;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_107;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_108;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_109;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_110;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_111;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_112;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_113;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_114;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_115;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_116;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_117;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_118;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_119;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_120;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_121;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_122;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_123;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_124;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_125;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_126;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_127;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_128;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_129;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_130;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_131;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_132;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_133;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_134;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_135;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_136;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_137;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_138;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_139;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_140;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_141;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_142;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_143;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_144;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_145;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_146;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_147;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_148;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_149;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_150;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_151;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_152;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_153;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_154;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_155;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_156;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_157;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_158;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_159;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_160;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_161;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_162;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_163;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_164;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_165;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_166;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_167;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_168;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_169;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_170;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_171;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_172;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_173;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_174;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_175;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_176;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_177;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_178;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_179;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_180;
  reg [31:0] bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_181;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_19;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_20;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_21;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_22;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_23;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_24;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_25;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_26;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_27;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_28;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_29;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_30;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_31;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_32;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_33;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_34;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_35;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_36;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_37;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_38;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_39;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_40;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_41;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_42;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_43;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_44;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_45;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_46;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_47;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_48;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_49;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_50;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_51;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_52;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_53;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_54;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_55;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_56;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_57;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_58;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_59;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_60;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_61;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_62;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_63;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_64;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_65;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_66;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_67;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_68;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_69;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_70;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_71;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_72;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_73;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_74;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_75;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_76;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_77;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_78;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_79;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_80;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_81;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_82;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_83;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_84;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_85;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_86;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_87;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_88;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_89;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_90;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_91;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_92;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_93;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_94;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_95;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_96;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_97;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_98;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_99;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_100;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_101;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_102;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_103;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_104;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_105;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_106;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_107;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_108;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_109;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_110;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_111;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_112;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_113;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_114;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_115;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_116;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_117;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_118;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_119;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_120;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_121;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_122;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_123;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_124;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_125;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_126;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_127;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_128;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_129;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_130;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_131;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_132;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_133;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_134;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_135;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_136;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_137;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_138;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_139;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_140;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_141;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_142;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_143;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_144;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_145;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_146;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_147;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_148;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_149;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_150;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_151;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_152;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_153;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_154;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_155;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_156;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_157;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_158;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_159;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_160;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_161;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_162;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_163;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_164;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_165;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_166;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_167;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_168;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_169;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_170;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_171;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_172;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_173;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_174;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_175;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_176;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_177;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_178;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_179;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_180;
  reg [31:0] dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_181;
  reg [31:0] bright_gauss_blur_1_update_0_stage_21;
  reg [31:0] bright_gauss_blur_1_update_0_stage_22;
  reg [31:0] bright_gauss_blur_1_update_0_stage_23;
  reg [31:0] bright_gauss_blur_1_update_0_stage_24;
  reg [31:0] bright_gauss_blur_1_update_0_stage_25;
  reg [31:0] bright_gauss_blur_1_update_0_stage_26;
  reg [31:0] bright_gauss_blur_1_update_0_stage_27;
  reg [31:0] bright_gauss_blur_1_update_0_stage_28;
  reg [31:0] bright_gauss_blur_1_update_0_stage_29;
  reg [31:0] bright_gauss_blur_1_update_0_stage_30;
  reg [31:0] bright_gauss_blur_1_update_0_stage_31;
  reg [31:0] bright_gauss_blur_1_update_0_stage_32;
  reg [31:0] bright_gauss_blur_1_update_0_stage_33;
  reg [31:0] bright_gauss_blur_1_update_0_stage_34;
  reg [31:0] bright_gauss_blur_1_update_0_stage_35;
  reg [31:0] bright_gauss_blur_1_update_0_stage_36;
  reg [31:0] bright_gauss_blur_1_update_0_stage_37;
  reg [31:0] bright_gauss_blur_1_update_0_stage_38;
  reg [31:0] bright_gauss_blur_1_update_0_stage_39;
  reg [31:0] bright_gauss_blur_1_update_0_stage_40;
  reg [31:0] bright_gauss_blur_1_update_0_stage_41;
  reg [31:0] bright_gauss_blur_1_update_0_stage_42;
  reg [31:0] bright_gauss_blur_1_update_0_stage_43;
  reg [31:0] bright_gauss_blur_1_update_0_stage_44;
  reg [31:0] bright_gauss_blur_1_update_0_stage_45;
  reg [31:0] bright_gauss_blur_1_update_0_stage_46;
  reg [31:0] bright_gauss_blur_1_update_0_stage_47;
  reg [31:0] bright_gauss_blur_1_update_0_stage_48;
  reg [31:0] bright_gauss_blur_1_update_0_stage_49;
  reg [31:0] bright_gauss_blur_1_update_0_stage_50;
  reg [31:0] bright_gauss_blur_1_update_0_stage_51;
  reg [31:0] bright_gauss_blur_1_update_0_stage_52;
  reg [31:0] bright_gauss_blur_1_update_0_stage_53;
  reg [31:0] bright_gauss_blur_1_update_0_stage_54;
  reg [31:0] bright_gauss_blur_1_update_0_stage_55;
  reg [31:0] bright_gauss_blur_1_update_0_stage_56;
  reg [31:0] bright_gauss_blur_1_update_0_stage_57;
  reg [31:0] bright_gauss_blur_1_update_0_stage_58;
  reg [31:0] bright_gauss_blur_1_update_0_stage_59;
  reg [31:0] bright_gauss_blur_1_update_0_stage_60;
  reg [31:0] bright_gauss_blur_1_update_0_stage_61;
  reg [31:0] bright_gauss_blur_1_update_0_stage_62;
  reg [31:0] bright_gauss_blur_1_update_0_stage_63;
  reg [31:0] bright_gauss_blur_1_update_0_stage_64;
  reg [31:0] bright_gauss_blur_1_update_0_stage_65;
  reg [31:0] bright_gauss_blur_1_update_0_stage_66;
  reg [31:0] bright_gauss_blur_1_update_0_stage_67;
  reg [31:0] bright_gauss_blur_1_update_0_stage_68;
  reg [31:0] bright_gauss_blur_1_update_0_stage_69;
  reg [31:0] bright_gauss_blur_1_update_0_stage_70;
  reg [31:0] bright_gauss_blur_1_update_0_stage_71;
  reg [31:0] bright_gauss_blur_1_update_0_stage_72;
  reg [31:0] bright_gauss_blur_1_update_0_stage_73;
  reg [31:0] bright_gauss_blur_1_update_0_stage_74;
  reg [31:0] bright_gauss_blur_1_update_0_stage_75;
  reg [31:0] bright_gauss_blur_1_update_0_stage_76;
  reg [31:0] bright_gauss_blur_1_update_0_stage_77;
  reg [31:0] bright_gauss_blur_1_update_0_stage_78;
  reg [31:0] bright_gauss_blur_1_update_0_stage_79;
  reg [31:0] bright_gauss_blur_1_update_0_stage_80;
  reg [31:0] bright_gauss_blur_1_update_0_stage_81;
  reg [31:0] bright_gauss_blur_1_update_0_stage_82;
  reg [31:0] bright_gauss_blur_1_update_0_stage_83;
  reg [31:0] bright_gauss_blur_1_update_0_stage_84;
  reg [31:0] bright_gauss_blur_1_update_0_stage_85;
  reg [31:0] bright_gauss_blur_1_update_0_stage_86;
  reg [31:0] bright_gauss_blur_1_update_0_stage_87;
  reg [31:0] bright_gauss_blur_1_update_0_stage_88;
  reg [31:0] bright_gauss_blur_1_update_0_stage_89;
  reg [31:0] bright_gauss_blur_1_update_0_stage_90;
  reg [31:0] bright_gauss_blur_1_update_0_stage_91;
  reg [31:0] bright_gauss_blur_1_update_0_stage_92;
  reg [31:0] bright_gauss_blur_1_update_0_stage_93;
  reg [31:0] bright_gauss_blur_1_update_0_stage_94;
  reg [31:0] bright_gauss_blur_1_update_0_stage_95;
  reg [31:0] bright_gauss_blur_1_update_0_stage_96;
  reg [31:0] bright_gauss_blur_1_update_0_stage_97;
  reg [31:0] bright_gauss_blur_1_update_0_stage_98;
  reg [31:0] bright_gauss_blur_1_update_0_stage_99;
  reg [31:0] bright_gauss_blur_1_update_0_stage_100;
  reg [31:0] bright_gauss_blur_1_update_0_stage_101;
  reg [31:0] bright_gauss_blur_1_update_0_stage_102;
  reg [31:0] bright_gauss_blur_1_update_0_stage_103;
  reg [31:0] bright_gauss_blur_1_update_0_stage_104;
  reg [31:0] bright_gauss_blur_1_update_0_stage_105;
  reg [31:0] bright_gauss_blur_1_update_0_stage_106;
  reg [31:0] bright_gauss_blur_1_update_0_stage_107;
  reg [31:0] bright_gauss_blur_1_update_0_stage_108;
  reg [31:0] bright_gauss_blur_1_update_0_stage_109;
  reg [31:0] bright_gauss_blur_1_update_0_stage_110;
  reg [31:0] bright_gauss_blur_1_update_0_stage_111;
  reg [31:0] bright_gauss_blur_1_update_0_stage_112;
  reg [31:0] bright_gauss_blur_1_update_0_stage_113;
  reg [31:0] bright_gauss_blur_1_update_0_stage_114;
  reg [31:0] bright_gauss_blur_1_update_0_stage_115;
  reg [31:0] bright_gauss_blur_1_update_0_stage_116;
  reg [31:0] bright_gauss_blur_1_update_0_stage_117;
  reg [31:0] bright_gauss_blur_1_update_0_stage_118;
  reg [31:0] bright_gauss_blur_1_update_0_stage_119;
  reg [31:0] bright_gauss_blur_1_update_0_stage_120;
  reg [31:0] bright_gauss_blur_1_update_0_stage_121;
  reg [31:0] bright_gauss_blur_1_update_0_stage_122;
  reg [31:0] bright_gauss_blur_1_update_0_stage_123;
  reg [31:0] bright_gauss_blur_1_update_0_stage_124;
  reg [31:0] bright_gauss_blur_1_update_0_stage_125;
  reg [31:0] bright_gauss_blur_1_update_0_stage_126;
  reg [31:0] bright_gauss_blur_1_update_0_stage_127;
  reg [31:0] bright_gauss_blur_1_update_0_stage_128;
  reg [31:0] bright_gauss_blur_1_update_0_stage_129;
  reg [31:0] bright_gauss_blur_1_update_0_stage_130;
  reg [31:0] bright_gauss_blur_1_update_0_stage_131;
  reg [31:0] bright_gauss_blur_1_update_0_stage_132;
  reg [31:0] bright_gauss_blur_1_update_0_stage_133;
  reg [31:0] bright_gauss_blur_1_update_0_stage_134;
  reg [31:0] bright_gauss_blur_1_update_0_stage_135;
  reg [31:0] bright_gauss_blur_1_update_0_stage_136;
  reg [31:0] bright_gauss_blur_1_update_0_stage_137;
  reg [31:0] bright_gauss_blur_1_update_0_stage_138;
  reg [31:0] bright_gauss_blur_1_update_0_stage_139;
  reg [31:0] bright_gauss_blur_1_update_0_stage_140;
  reg [31:0] bright_gauss_blur_1_update_0_stage_141;
  reg [31:0] bright_gauss_blur_1_update_0_stage_142;
  reg [31:0] bright_gauss_blur_1_update_0_stage_143;
  reg [31:0] bright_gauss_blur_1_update_0_stage_144;
  reg [31:0] bright_gauss_blur_1_update_0_stage_145;
  reg [31:0] bright_gauss_blur_1_update_0_stage_146;
  reg [31:0] bright_gauss_blur_1_update_0_stage_147;
  reg [31:0] bright_gauss_blur_1_update_0_stage_148;
  reg [31:0] bright_gauss_blur_1_update_0_stage_149;
  reg [31:0] bright_gauss_blur_1_update_0_stage_150;
  reg [31:0] bright_gauss_blur_1_update_0_stage_151;
  reg [31:0] bright_gauss_blur_1_update_0_stage_152;
  reg [31:0] bright_gauss_blur_1_update_0_stage_153;
  reg [31:0] bright_gauss_blur_1_update_0_stage_154;
  reg [31:0] bright_gauss_blur_1_update_0_stage_155;
  reg [31:0] bright_gauss_blur_1_update_0_stage_156;
  reg [31:0] bright_gauss_blur_1_update_0_stage_157;
  reg [31:0] bright_gauss_blur_1_update_0_stage_158;
  reg [31:0] bright_gauss_blur_1_update_0_stage_159;
  reg [31:0] bright_gauss_blur_1_update_0_stage_160;
  reg [31:0] bright_gauss_blur_1_update_0_stage_161;
  reg [31:0] bright_gauss_blur_1_update_0_stage_162;
  reg [31:0] bright_gauss_blur_1_update_0_stage_163;
  reg [31:0] bright_gauss_blur_1_update_0_stage_164;
  reg [31:0] bright_gauss_blur_1_update_0_stage_165;
  reg [31:0] bright_gauss_blur_1_update_0_stage_166;
  reg [31:0] bright_gauss_blur_1_update_0_stage_167;
  reg [31:0] bright_gauss_blur_1_update_0_stage_168;
  reg [31:0] bright_gauss_blur_1_update_0_stage_169;
  reg [31:0] bright_gauss_blur_1_update_0_stage_170;
  reg [31:0] bright_gauss_blur_1_update_0_stage_171;
  reg [31:0] bright_gauss_blur_1_update_0_stage_172;
  reg [31:0] bright_gauss_blur_1_update_0_stage_173;
  reg [31:0] bright_gauss_blur_1_update_0_stage_174;
  reg [31:0] bright_gauss_blur_1_update_0_stage_175;
  reg [31:0] bright_gauss_blur_1_update_0_stage_176;
  reg [31:0] bright_gauss_blur_1_update_0_stage_177;
  reg [31:0] bright_gauss_blur_1_update_0_stage_178;
  reg [31:0] bright_gauss_blur_1_update_0_stage_179;
  reg [31:0] bright_gauss_blur_1_update_0_stage_180;
  reg [31:0] bright_gauss_blur_1_update_0_stage_181;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_20;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_21;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_22;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_23;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_24;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_25;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_26;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_27;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_28;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_29;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_30;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_31;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_32;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_33;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_34;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_35;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_36;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_37;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_38;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_39;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_40;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_41;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_42;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_43;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_44;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_45;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_46;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_47;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_48;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_49;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_50;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_51;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_52;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_53;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_54;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_55;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_56;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_57;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_58;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_59;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_60;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_61;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_62;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_63;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_64;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_65;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_66;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_67;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_68;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_69;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_70;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_71;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_72;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_73;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_74;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_75;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_76;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_77;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_78;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_79;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_80;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_81;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_82;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_83;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_84;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_85;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_86;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_87;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_88;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_89;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_90;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_91;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_92;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_93;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_94;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_95;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_96;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_97;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_98;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_99;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_100;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_101;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_102;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_103;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_104;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_105;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_106;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_107;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_108;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_109;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_110;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_111;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_112;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_113;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_114;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_115;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_116;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_117;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_118;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_119;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_120;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_121;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_122;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_123;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_124;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_125;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_126;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_127;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_128;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_129;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_130;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_131;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_132;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_133;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_134;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_135;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_136;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_137;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_138;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_139;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_140;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_141;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_142;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_143;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_144;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_145;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_146;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_147;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_148;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_149;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_150;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_151;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_152;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_153;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_154;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_155;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_156;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_157;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_158;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_159;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_160;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_161;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_162;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_163;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_164;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_165;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_166;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_167;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_168;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_169;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_170;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_171;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_172;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_173;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_174;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_175;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_176;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_177;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_178;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_179;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_180;
  reg [287:0] bright_bright_gauss_blur_1_update_0_read_read_12_stage_181;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_22;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_23;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_24;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_25;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_26;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_27;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_28;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_29;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_30;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_31;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_32;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_33;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_34;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_35;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_36;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_37;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_38;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_39;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_40;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_41;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_42;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_43;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_44;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_45;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_46;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_47;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_48;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_49;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_50;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_51;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_52;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_53;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_54;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_55;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_56;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_57;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_58;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_59;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_60;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_61;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_62;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_63;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_64;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_65;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_66;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_67;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_68;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_69;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_70;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_71;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_72;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_73;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_74;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_75;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_76;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_77;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_78;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_79;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_80;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_81;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_82;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_83;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_84;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_85;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_86;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_87;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_88;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_89;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_90;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_91;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_92;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_93;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_94;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_95;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_96;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_97;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_98;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_99;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_100;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_101;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_102;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_103;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_104;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_105;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_106;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_107;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_108;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_109;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_110;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_111;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_112;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_113;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_114;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_115;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_116;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_117;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_118;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_119;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_120;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_121;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_122;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_123;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_124;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_125;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_126;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_127;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_128;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_129;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_130;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_131;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_132;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_133;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_134;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_135;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_136;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_137;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_138;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_139;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_140;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_141;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_142;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_143;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_144;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_145;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_146;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_147;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_148;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_149;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_150;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_151;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_152;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_153;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_154;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_155;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_156;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_157;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_158;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_159;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_160;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_161;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_162;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_163;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_164;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_165;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_166;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_167;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_168;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_169;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_170;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_171;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_172;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_173;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_174;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_175;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_176;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_177;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_178;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_179;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_180;
  reg [31:0] bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_181;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_61;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_62;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_63;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_64;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_65;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_66;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_67;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_68;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_69;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_70;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_71;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_72;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_73;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_74;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_75;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_76;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_77;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_78;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_79;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_80;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_81;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_82;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_83;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_84;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_85;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_86;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_87;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_88;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_89;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_90;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_91;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_92;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_93;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_94;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_95;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_96;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_97;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_98;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_99;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_100;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_101;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_102;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_103;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_104;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_105;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_106;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_107;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_108;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_109;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_110;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_111;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_112;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_113;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_114;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_115;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_116;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_117;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_118;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_119;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_120;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_121;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_122;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_123;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_124;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_125;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_126;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_127;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_128;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_129;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_130;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_131;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_132;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_133;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_134;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_135;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_136;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_137;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_138;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_139;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_140;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_141;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_142;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_143;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_144;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_145;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_146;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_147;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_148;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_149;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_150;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_151;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_152;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_153;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_154;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_155;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_156;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_157;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_158;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_159;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_160;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_161;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_162;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_163;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_164;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_165;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_166;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_167;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_168;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_169;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_170;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_171;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_172;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_173;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_174;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_175;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_176;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_177;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_178;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_179;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_180;
  reg [31:0] bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_181;
  reg [31:0] bright_laplace_us_1_update_0_stage_62;
  reg [31:0] bright_laplace_us_1_update_0_stage_63;
  reg [31:0] bright_laplace_us_1_update_0_stage_64;
  reg [31:0] bright_laplace_us_1_update_0_stage_65;
  reg [31:0] bright_laplace_us_1_update_0_stage_66;
  reg [31:0] bright_laplace_us_1_update_0_stage_67;
  reg [31:0] bright_laplace_us_1_update_0_stage_68;
  reg [31:0] bright_laplace_us_1_update_0_stage_69;
  reg [31:0] bright_laplace_us_1_update_0_stage_70;
  reg [31:0] bright_laplace_us_1_update_0_stage_71;
  reg [31:0] bright_laplace_us_1_update_0_stage_72;
  reg [31:0] bright_laplace_us_1_update_0_stage_73;
  reg [31:0] bright_laplace_us_1_update_0_stage_74;
  reg [31:0] bright_laplace_us_1_update_0_stage_75;
  reg [31:0] bright_laplace_us_1_update_0_stage_76;
  reg [31:0] bright_laplace_us_1_update_0_stage_77;
  reg [31:0] bright_laplace_us_1_update_0_stage_78;
  reg [31:0] bright_laplace_us_1_update_0_stage_79;
  reg [31:0] bright_laplace_us_1_update_0_stage_80;
  reg [31:0] bright_laplace_us_1_update_0_stage_81;
  reg [31:0] bright_laplace_us_1_update_0_stage_82;
  reg [31:0] bright_laplace_us_1_update_0_stage_83;
  reg [31:0] bright_laplace_us_1_update_0_stage_84;
  reg [31:0] bright_laplace_us_1_update_0_stage_85;
  reg [31:0] bright_laplace_us_1_update_0_stage_86;
  reg [31:0] bright_laplace_us_1_update_0_stage_87;
  reg [31:0] bright_laplace_us_1_update_0_stage_88;
  reg [31:0] bright_laplace_us_1_update_0_stage_89;
  reg [31:0] bright_laplace_us_1_update_0_stage_90;
  reg [31:0] bright_laplace_us_1_update_0_stage_91;
  reg [31:0] bright_laplace_us_1_update_0_stage_92;
  reg [31:0] bright_laplace_us_1_update_0_stage_93;
  reg [31:0] bright_laplace_us_1_update_0_stage_94;
  reg [31:0] bright_laplace_us_1_update_0_stage_95;
  reg [31:0] bright_laplace_us_1_update_0_stage_96;
  reg [31:0] bright_laplace_us_1_update_0_stage_97;
  reg [31:0] bright_laplace_us_1_update_0_stage_98;
  reg [31:0] bright_laplace_us_1_update_0_stage_99;
  reg [31:0] bright_laplace_us_1_update_0_stage_100;
  reg [31:0] bright_laplace_us_1_update_0_stage_101;
  reg [31:0] bright_laplace_us_1_update_0_stage_102;
  reg [31:0] bright_laplace_us_1_update_0_stage_103;
  reg [31:0] bright_laplace_us_1_update_0_stage_104;
  reg [31:0] bright_laplace_us_1_update_0_stage_105;
  reg [31:0] bright_laplace_us_1_update_0_stage_106;
  reg [31:0] bright_laplace_us_1_update_0_stage_107;
  reg [31:0] bright_laplace_us_1_update_0_stage_108;
  reg [31:0] bright_laplace_us_1_update_0_stage_109;
  reg [31:0] bright_laplace_us_1_update_0_stage_110;
  reg [31:0] bright_laplace_us_1_update_0_stage_111;
  reg [31:0] bright_laplace_us_1_update_0_stage_112;
  reg [31:0] bright_laplace_us_1_update_0_stage_113;
  reg [31:0] bright_laplace_us_1_update_0_stage_114;
  reg [31:0] bright_laplace_us_1_update_0_stage_115;
  reg [31:0] bright_laplace_us_1_update_0_stage_116;
  reg [31:0] bright_laplace_us_1_update_0_stage_117;
  reg [31:0] bright_laplace_us_1_update_0_stage_118;
  reg [31:0] bright_laplace_us_1_update_0_stage_119;
  reg [31:0] bright_laplace_us_1_update_0_stage_120;
  reg [31:0] bright_laplace_us_1_update_0_stage_121;
  reg [31:0] bright_laplace_us_1_update_0_stage_122;
  reg [31:0] bright_laplace_us_1_update_0_stage_123;
  reg [31:0] bright_laplace_us_1_update_0_stage_124;
  reg [31:0] bright_laplace_us_1_update_0_stage_125;
  reg [31:0] bright_laplace_us_1_update_0_stage_126;
  reg [31:0] bright_laplace_us_1_update_0_stage_127;
  reg [31:0] bright_laplace_us_1_update_0_stage_128;
  reg [31:0] bright_laplace_us_1_update_0_stage_129;
  reg [31:0] bright_laplace_us_1_update_0_stage_130;
  reg [31:0] bright_laplace_us_1_update_0_stage_131;
  reg [31:0] bright_laplace_us_1_update_0_stage_132;
  reg [31:0] bright_laplace_us_1_update_0_stage_133;
  reg [31:0] bright_laplace_us_1_update_0_stage_134;
  reg [31:0] bright_laplace_us_1_update_0_stage_135;
  reg [31:0] bright_laplace_us_1_update_0_stage_136;
  reg [31:0] bright_laplace_us_1_update_0_stage_137;
  reg [31:0] bright_laplace_us_1_update_0_stage_138;
  reg [31:0] bright_laplace_us_1_update_0_stage_139;
  reg [31:0] bright_laplace_us_1_update_0_stage_140;
  reg [31:0] bright_laplace_us_1_update_0_stage_141;
  reg [31:0] bright_laplace_us_1_update_0_stage_142;
  reg [31:0] bright_laplace_us_1_update_0_stage_143;
  reg [31:0] bright_laplace_us_1_update_0_stage_144;
  reg [31:0] bright_laplace_us_1_update_0_stage_145;
  reg [31:0] bright_laplace_us_1_update_0_stage_146;
  reg [31:0] bright_laplace_us_1_update_0_stage_147;
  reg [31:0] bright_laplace_us_1_update_0_stage_148;
  reg [31:0] bright_laplace_us_1_update_0_stage_149;
  reg [31:0] bright_laplace_us_1_update_0_stage_150;
  reg [31:0] bright_laplace_us_1_update_0_stage_151;
  reg [31:0] bright_laplace_us_1_update_0_stage_152;
  reg [31:0] bright_laplace_us_1_update_0_stage_153;
  reg [31:0] bright_laplace_us_1_update_0_stage_154;
  reg [31:0] bright_laplace_us_1_update_0_stage_155;
  reg [31:0] bright_laplace_us_1_update_0_stage_156;
  reg [31:0] bright_laplace_us_1_update_0_stage_157;
  reg [31:0] bright_laplace_us_1_update_0_stage_158;
  reg [31:0] bright_laplace_us_1_update_0_stage_159;
  reg [31:0] bright_laplace_us_1_update_0_stage_160;
  reg [31:0] bright_laplace_us_1_update_0_stage_161;
  reg [31:0] bright_laplace_us_1_update_0_stage_162;
  reg [31:0] bright_laplace_us_1_update_0_stage_163;
  reg [31:0] bright_laplace_us_1_update_0_stage_164;
  reg [31:0] bright_laplace_us_1_update_0_stage_165;
  reg [31:0] bright_laplace_us_1_update_0_stage_166;
  reg [31:0] bright_laplace_us_1_update_0_stage_167;
  reg [31:0] bright_laplace_us_1_update_0_stage_168;
  reg [31:0] bright_laplace_us_1_update_0_stage_169;
  reg [31:0] bright_laplace_us_1_update_0_stage_170;
  reg [31:0] bright_laplace_us_1_update_0_stage_171;
  reg [31:0] bright_laplace_us_1_update_0_stage_172;
  reg [31:0] bright_laplace_us_1_update_0_stage_173;
  reg [31:0] bright_laplace_us_1_update_0_stage_174;
  reg [31:0] bright_laplace_us_1_update_0_stage_175;
  reg [31:0] bright_laplace_us_1_update_0_stage_176;
  reg [31:0] bright_laplace_us_1_update_0_stage_177;
  reg [31:0] bright_laplace_us_1_update_0_stage_178;
  reg [31:0] bright_laplace_us_1_update_0_stage_179;
  reg [31:0] bright_laplace_us_1_update_0_stage_180;
  reg [31:0] bright_laplace_us_1_update_0_stage_181;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_63;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_64;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_65;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_66;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_67;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_68;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_69;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_70;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_71;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_72;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_73;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_74;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_75;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_76;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_77;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_78;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_79;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_80;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_81;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_82;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_83;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_84;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_85;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_86;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_87;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_88;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_89;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_90;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_91;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_92;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_93;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_94;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_95;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_96;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_97;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_98;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_99;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_100;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_101;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_102;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_103;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_104;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_105;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_106;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_107;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_108;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_109;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_110;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_111;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_112;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_113;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_114;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_115;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_116;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_117;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_118;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_119;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_120;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_121;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_122;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_123;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_124;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_125;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_126;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_127;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_128;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_129;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_130;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_131;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_132;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_133;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_134;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_135;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_136;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_137;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_138;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_139;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_140;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_141;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_142;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_143;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_144;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_145;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_146;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_147;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_148;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_149;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_150;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_151;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_152;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_153;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_154;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_155;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_156;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_157;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_158;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_159;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_160;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_161;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_162;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_163;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_164;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_165;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_166;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_167;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_168;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_169;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_170;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_171;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_172;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_173;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_174;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_175;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_176;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_177;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_178;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_179;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_180;
  reg [31:0] bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_83;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_84;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_85;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_86;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_87;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_88;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_89;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_90;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_91;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_92;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_93;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_94;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_95;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_96;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_97;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_98;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_99;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_100;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_101;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_102;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_103;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_104;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_105;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_106;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_107;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_108;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_109;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_110;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_111;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_112;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_113;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_114;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_115;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_116;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_117;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_118;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_119;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_120;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_121;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_122;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_123;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_124;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_125;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_126;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_127;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_128;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_129;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_130;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_131;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_132;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_133;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_134;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_135;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_136;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_137;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_138;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_1_update_0_stage_181;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_82;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_83;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_84;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_85;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_86;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_87;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_88;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_89;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_90;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_91;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_92;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_93;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_94;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_95;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_96;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_97;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_98;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_99;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_100;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_101;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_102;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_103;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_104;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_105;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_106;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_107;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_108;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_109;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_110;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_111;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_112;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_113;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_114;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_115;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_116;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_117;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_118;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_119;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_120;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_121;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_122;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_123;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_124;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_125;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_126;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_127;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_128;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_129;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_130;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_131;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_132;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_133;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_134;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_135;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_136;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_137;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_138;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_139;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_140;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_141;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_142;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_143;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_144;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_145;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_146;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_147;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_148;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_149;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_150;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_151;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_152;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_153;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_154;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_155;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_156;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_157;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_158;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_159;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_160;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_161;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_162;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_163;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_164;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_165;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_166;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_167;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_168;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_169;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_170;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_171;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_172;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_173;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_174;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_175;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_176;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_177;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_178;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_179;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_180;
  reg [287:0] bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_181;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_88;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_89;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_90;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_91;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_92;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_93;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_94;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_95;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_96;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_97;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_98;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_99;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_100;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_101;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_102;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_103;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_104;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_105;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_106;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_107;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_108;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_109;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_110;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_111;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_112;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_113;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_114;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_115;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_116;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_117;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_118;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_119;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_120;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_121;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_122;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_123;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_124;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_125;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_126;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_127;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_128;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_129;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_130;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_131;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_132;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_133;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_134;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_135;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_136;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_137;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_138;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_139;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_140;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_141;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_142;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_143;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_144;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_145;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_146;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_147;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_148;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_149;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_150;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_151;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_152;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_153;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_154;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_155;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_156;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_157;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_158;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_159;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_160;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_161;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_162;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_163;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_164;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_165;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_166;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_167;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_168;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_169;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_170;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_171;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_172;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_173;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_174;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_175;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_176;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_177;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_178;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_179;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_180;
  reg [31:0] bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_84;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_85;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_86;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_87;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_88;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_89;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_90;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_91;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_92;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_93;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_94;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_95;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_96;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_97;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_98;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_99;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_100;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_101;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_102;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_103;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_104;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_105;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_106;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_107;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_108;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_109;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_110;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_111;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_112;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_113;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_114;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_115;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_116;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_117;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_118;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_119;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_120;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_121;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_122;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_123;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_124;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_125;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_126;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_127;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_128;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_129;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_130;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_131;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_132;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_133;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_134;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_135;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_136;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_137;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_138;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_181;
  reg [31:0] bright_laplace_us_2_update_0_stage_89;
  reg [31:0] bright_laplace_us_2_update_0_stage_90;
  reg [31:0] bright_laplace_us_2_update_0_stage_91;
  reg [31:0] bright_laplace_us_2_update_0_stage_92;
  reg [31:0] bright_laplace_us_2_update_0_stage_93;
  reg [31:0] bright_laplace_us_2_update_0_stage_94;
  reg [31:0] bright_laplace_us_2_update_0_stage_95;
  reg [31:0] bright_laplace_us_2_update_0_stage_96;
  reg [31:0] bright_laplace_us_2_update_0_stage_97;
  reg [31:0] bright_laplace_us_2_update_0_stage_98;
  reg [31:0] bright_laplace_us_2_update_0_stage_99;
  reg [31:0] bright_laplace_us_2_update_0_stage_100;
  reg [31:0] bright_laplace_us_2_update_0_stage_101;
  reg [31:0] bright_laplace_us_2_update_0_stage_102;
  reg [31:0] bright_laplace_us_2_update_0_stage_103;
  reg [31:0] bright_laplace_us_2_update_0_stage_104;
  reg [31:0] bright_laplace_us_2_update_0_stage_105;
  reg [31:0] bright_laplace_us_2_update_0_stage_106;
  reg [31:0] bright_laplace_us_2_update_0_stage_107;
  reg [31:0] bright_laplace_us_2_update_0_stage_108;
  reg [31:0] bright_laplace_us_2_update_0_stage_109;
  reg [31:0] bright_laplace_us_2_update_0_stage_110;
  reg [31:0] bright_laplace_us_2_update_0_stage_111;
  reg [31:0] bright_laplace_us_2_update_0_stage_112;
  reg [31:0] bright_laplace_us_2_update_0_stage_113;
  reg [31:0] bright_laplace_us_2_update_0_stage_114;
  reg [31:0] bright_laplace_us_2_update_0_stage_115;
  reg [31:0] bright_laplace_us_2_update_0_stage_116;
  reg [31:0] bright_laplace_us_2_update_0_stage_117;
  reg [31:0] bright_laplace_us_2_update_0_stage_118;
  reg [31:0] bright_laplace_us_2_update_0_stage_119;
  reg [31:0] bright_laplace_us_2_update_0_stage_120;
  reg [31:0] bright_laplace_us_2_update_0_stage_121;
  reg [31:0] bright_laplace_us_2_update_0_stage_122;
  reg [31:0] bright_laplace_us_2_update_0_stage_123;
  reg [31:0] bright_laplace_us_2_update_0_stage_124;
  reg [31:0] bright_laplace_us_2_update_0_stage_125;
  reg [31:0] bright_laplace_us_2_update_0_stage_126;
  reg [31:0] bright_laplace_us_2_update_0_stage_127;
  reg [31:0] bright_laplace_us_2_update_0_stage_128;
  reg [31:0] bright_laplace_us_2_update_0_stage_129;
  reg [31:0] bright_laplace_us_2_update_0_stage_130;
  reg [31:0] bright_laplace_us_2_update_0_stage_131;
  reg [31:0] bright_laplace_us_2_update_0_stage_132;
  reg [31:0] bright_laplace_us_2_update_0_stage_133;
  reg [31:0] bright_laplace_us_2_update_0_stage_134;
  reg [31:0] bright_laplace_us_2_update_0_stage_135;
  reg [31:0] bright_laplace_us_2_update_0_stage_136;
  reg [31:0] bright_laplace_us_2_update_0_stage_137;
  reg [31:0] bright_laplace_us_2_update_0_stage_138;
  reg [31:0] bright_laplace_us_2_update_0_stage_139;
  reg [31:0] bright_laplace_us_2_update_0_stage_140;
  reg [31:0] bright_laplace_us_2_update_0_stage_141;
  reg [31:0] bright_laplace_us_2_update_0_stage_142;
  reg [31:0] bright_laplace_us_2_update_0_stage_143;
  reg [31:0] bright_laplace_us_2_update_0_stage_144;
  reg [31:0] bright_laplace_us_2_update_0_stage_145;
  reg [31:0] bright_laplace_us_2_update_0_stage_146;
  reg [31:0] bright_laplace_us_2_update_0_stage_147;
  reg [31:0] bright_laplace_us_2_update_0_stage_148;
  reg [31:0] bright_laplace_us_2_update_0_stage_149;
  reg [31:0] bright_laplace_us_2_update_0_stage_150;
  reg [31:0] bright_laplace_us_2_update_0_stage_151;
  reg [31:0] bright_laplace_us_2_update_0_stage_152;
  reg [31:0] bright_laplace_us_2_update_0_stage_153;
  reg [31:0] bright_laplace_us_2_update_0_stage_154;
  reg [31:0] bright_laplace_us_2_update_0_stage_155;
  reg [31:0] bright_laplace_us_2_update_0_stage_156;
  reg [31:0] bright_laplace_us_2_update_0_stage_157;
  reg [31:0] bright_laplace_us_2_update_0_stage_158;
  reg [31:0] bright_laplace_us_2_update_0_stage_159;
  reg [31:0] bright_laplace_us_2_update_0_stage_160;
  reg [31:0] bright_laplace_us_2_update_0_stage_161;
  reg [31:0] bright_laplace_us_2_update_0_stage_162;
  reg [31:0] bright_laplace_us_2_update_0_stage_163;
  reg [31:0] bright_laplace_us_2_update_0_stage_164;
  reg [31:0] bright_laplace_us_2_update_0_stage_165;
  reg [31:0] bright_laplace_us_2_update_0_stage_166;
  reg [31:0] bright_laplace_us_2_update_0_stage_167;
  reg [31:0] bright_laplace_us_2_update_0_stage_168;
  reg [31:0] bright_laplace_us_2_update_0_stage_169;
  reg [31:0] bright_laplace_us_2_update_0_stage_170;
  reg [31:0] bright_laplace_us_2_update_0_stage_171;
  reg [31:0] bright_laplace_us_2_update_0_stage_172;
  reg [31:0] bright_laplace_us_2_update_0_stage_173;
  reg [31:0] bright_laplace_us_2_update_0_stage_174;
  reg [31:0] bright_laplace_us_2_update_0_stage_175;
  reg [31:0] bright_laplace_us_2_update_0_stage_176;
  reg [31:0] bright_laplace_us_2_update_0_stage_177;
  reg [31:0] bright_laplace_us_2_update_0_stage_178;
  reg [31:0] bright_laplace_us_2_update_0_stage_179;
  reg [31:0] bright_laplace_us_2_update_0_stage_180;
  reg [31:0] bright_laplace_us_2_update_0_stage_181;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_90;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_91;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_92;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_93;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_94;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_95;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_96;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_97;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_98;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_99;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_100;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_101;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_102;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_103;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_104;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_105;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_106;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_107;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_108;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_109;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_110;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_111;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_112;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_113;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_114;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_115;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_116;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_117;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_118;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_119;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_120;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_121;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_122;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_123;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_124;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_125;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_126;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_127;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_128;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_129;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_130;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_131;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_132;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_133;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_134;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_135;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_136;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_137;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_138;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_139;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_140;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_141;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_142;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_143;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_144;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_145;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_146;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_147;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_148;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_149;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_150;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_151;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_152;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_153;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_154;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_155;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_156;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_157;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_158;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_159;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_160;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_161;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_162;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_163;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_164;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_165;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_166;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_167;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_168;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_169;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_170;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_171;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_172;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_173;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_174;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_175;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_176;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_177;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_178;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_179;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_180;
  reg [31:0] bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_181;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_91;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_92;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_93;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_94;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_95;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_96;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_97;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_98;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_99;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_100;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_101;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_102;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_103;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_104;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_105;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_106;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_107;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_108;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_109;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_110;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_111;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_112;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_113;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_114;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_115;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_116;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_117;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_118;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_119;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_120;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_121;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_122;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_123;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_124;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_125;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_126;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_127;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_128;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_129;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_130;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_131;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_132;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_133;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_134;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_135;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_136;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_137;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_138;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_139;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_140;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_141;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_142;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_143;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_144;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_145;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_146;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_147;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_148;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_149;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_150;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_151;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_152;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_153;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_154;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_155;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_156;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_157;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_158;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_159;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_160;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_161;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_162;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_163;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_164;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_165;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_166;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_167;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_168;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_169;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_170;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_171;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_172;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_173;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_174;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_175;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_176;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_177;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_178;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_179;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_180;
  reg [31:0] dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_181;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_148;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_149;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_150;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_151;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_152;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_153;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_154;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_155;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_156;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_157;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_158;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_159;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_160;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_161;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_162;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_163;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_164;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_165;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_166;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_167;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_168;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_169;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_170;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_171;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_172;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_173;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_174;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_175;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_176;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_177;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_178;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_179;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_180;
  reg [31:0] dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_181;
  reg [31:0] fused_level_3_update_0_stage_165;
  reg [31:0] fused_level_3_update_0_stage_166;
  reg [31:0] fused_level_3_update_0_stage_167;
  reg [31:0] fused_level_3_update_0_stage_168;
  reg [31:0] fused_level_3_update_0_stage_169;
  reg [31:0] fused_level_3_update_0_stage_170;
  reg [31:0] fused_level_3_update_0_stage_171;
  reg [31:0] fused_level_3_update_0_stage_172;
  reg [31:0] fused_level_3_update_0_stage_173;
  reg [31:0] fused_level_3_update_0_stage_174;
  reg [31:0] fused_level_3_update_0_stage_175;
  reg [31:0] fused_level_3_update_0_stage_176;
  reg [31:0] fused_level_3_update_0_stage_177;
  reg [31:0] fused_level_3_update_0_stage_178;
  reg [31:0] fused_level_3_update_0_stage_179;
  reg [31:0] fused_level_3_update_0_stage_180;
  reg [31:0] fused_level_3_update_0_stage_181;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_166;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_167;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_168;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_169;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_170;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_171;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_172;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_173;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_174;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_175;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_176;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_177;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_178;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_179;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_180;
  reg [31:0] fused_level_3_fused_level_3_update_0_write_write_116_stage_181;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_167;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_168;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_169;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_170;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_171;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_172;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_173;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_174;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_175;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_176;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_177;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_178;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_179;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_180;
  reg [31:0] fused_level_3_final_merged_2_update_0_read_read_117_stage_181;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_168;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_169;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_170;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_171;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_172;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_173;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_174;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_175;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_176;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_177;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_178;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_179;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_180;
  reg [31:0] fused_level_2_final_merged_2_update_0_read_read_118_stage_181;
  reg [31:0] final_merged_2_update_0_stage_169;
  reg [31:0] final_merged_2_update_0_stage_170;
  reg [31:0] final_merged_2_update_0_stage_171;
  reg [31:0] final_merged_2_update_0_stage_172;
  reg [31:0] final_merged_2_update_0_stage_173;
  reg [31:0] final_merged_2_update_0_stage_174;
  reg [31:0] final_merged_2_update_0_stage_175;
  reg [31:0] final_merged_2_update_0_stage_176;
  reg [31:0] final_merged_2_update_0_stage_177;
  reg [31:0] final_merged_2_update_0_stage_178;
  reg [31:0] final_merged_2_update_0_stage_179;
  reg [31:0] final_merged_2_update_0_stage_180;
  reg [31:0] final_merged_2_update_0_stage_181;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_170;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_171;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_172;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_173;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_174;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_175;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_176;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_177;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_178;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_179;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_180;
  reg [31:0] final_merged_2_final_merged_2_update_0_write_write_119_stage_181;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_175;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_176;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_177;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_178;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_179;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_180;
  reg [31:0] final_merged_1_final_merged_0_update_0_read_read_123_stage_181;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_176;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_177;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_178;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_179;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_180;
  reg [31:0] fused_level_0_final_merged_0_update_0_read_read_124_stage_181;
  reg [31:0] final_merged_0_update_0_stage_177;
  reg [31:0] final_merged_0_update_0_stage_178;
  reg [31:0] final_merged_0_update_0_stage_179;
  reg [31:0] final_merged_0_update_0_stage_180;
  reg [31:0] final_merged_0_update_0_stage_181;
  reg [31:0] final_merged_0_final_merged_0_update_0_write_write_125_stage_178;
  reg [31:0] final_merged_0_final_merged_0_update_0_write_write_125_stage_179;
  reg [31:0] final_merged_0_final_merged_0_update_0_write_write_125_stage_180;
  reg [31:0] final_merged_0_final_merged_0_update_0_write_write_125_stage_181;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_26;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_27;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_28;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_29;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_30;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_31;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_32;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_33;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_34;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_35;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_36;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_37;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_38;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_39;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_40;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_41;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_42;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_43;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_44;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_45;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_46;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_47;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_48;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_49;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_50;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_51;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_52;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_53;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_54;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_55;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_56;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_57;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_58;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_59;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_60;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_61;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_62;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_63;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_64;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_65;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_66;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_67;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_68;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_69;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_70;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_71;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_72;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_73;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_74;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_75;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_76;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_77;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_78;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_79;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_80;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_81;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_82;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_83;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_84;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_85;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_86;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_87;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_88;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_89;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_90;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_91;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_92;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_93;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_94;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_95;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_96;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_97;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_98;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_99;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_100;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_101;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_102;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_103;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_104;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_105;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_106;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_107;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_108;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_109;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_110;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_111;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_112;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_113;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_114;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_115;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_116;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_117;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_118;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_119;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_120;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_121;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_122;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_123;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_124;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_125;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_126;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_127;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_128;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_129;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_130;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_131;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_132;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_133;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_134;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_135;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_136;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_137;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_138;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_139;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_140;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_141;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_142;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_143;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_144;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_145;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_146;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_147;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_148;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_149;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_150;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_151;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_152;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_153;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_154;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_155;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_156;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_157;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_158;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_159;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_160;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_161;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_162;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_163;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_164;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_165;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_166;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_167;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_168;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_169;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_170;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_171;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_172;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_173;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_174;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_175;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_176;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_177;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_178;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_179;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_180;
  reg [31:0] dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_181;
  reg [31:0] dark_laplace_us_0_update_0_stage_27;
  reg [31:0] dark_laplace_us_0_update_0_stage_28;
  reg [31:0] dark_laplace_us_0_update_0_stage_29;
  reg [31:0] dark_laplace_us_0_update_0_stage_30;
  reg [31:0] dark_laplace_us_0_update_0_stage_31;
  reg [31:0] dark_laplace_us_0_update_0_stage_32;
  reg [31:0] dark_laplace_us_0_update_0_stage_33;
  reg [31:0] dark_laplace_us_0_update_0_stage_34;
  reg [31:0] dark_laplace_us_0_update_0_stage_35;
  reg [31:0] dark_laplace_us_0_update_0_stage_36;
  reg [31:0] dark_laplace_us_0_update_0_stage_37;
  reg [31:0] dark_laplace_us_0_update_0_stage_38;
  reg [31:0] dark_laplace_us_0_update_0_stage_39;
  reg [31:0] dark_laplace_us_0_update_0_stage_40;
  reg [31:0] dark_laplace_us_0_update_0_stage_41;
  reg [31:0] dark_laplace_us_0_update_0_stage_42;
  reg [31:0] dark_laplace_us_0_update_0_stage_43;
  reg [31:0] dark_laplace_us_0_update_0_stage_44;
  reg [31:0] dark_laplace_us_0_update_0_stage_45;
  reg [31:0] dark_laplace_us_0_update_0_stage_46;
  reg [31:0] dark_laplace_us_0_update_0_stage_47;
  reg [31:0] dark_laplace_us_0_update_0_stage_48;
  reg [31:0] dark_laplace_us_0_update_0_stage_49;
  reg [31:0] dark_laplace_us_0_update_0_stage_50;
  reg [31:0] dark_laplace_us_0_update_0_stage_51;
  reg [31:0] dark_laplace_us_0_update_0_stage_52;
  reg [31:0] dark_laplace_us_0_update_0_stage_53;
  reg [31:0] dark_laplace_us_0_update_0_stage_54;
  reg [31:0] dark_laplace_us_0_update_0_stage_55;
  reg [31:0] dark_laplace_us_0_update_0_stage_56;
  reg [31:0] dark_laplace_us_0_update_0_stage_57;
  reg [31:0] dark_laplace_us_0_update_0_stage_58;
  reg [31:0] dark_laplace_us_0_update_0_stage_59;
  reg [31:0] dark_laplace_us_0_update_0_stage_60;
  reg [31:0] dark_laplace_us_0_update_0_stage_61;
  reg [31:0] dark_laplace_us_0_update_0_stage_62;
  reg [31:0] dark_laplace_us_0_update_0_stage_63;
  reg [31:0] dark_laplace_us_0_update_0_stage_64;
  reg [31:0] dark_laplace_us_0_update_0_stage_65;
  reg [31:0] dark_laplace_us_0_update_0_stage_66;
  reg [31:0] dark_laplace_us_0_update_0_stage_67;
  reg [31:0] dark_laplace_us_0_update_0_stage_68;
  reg [31:0] dark_laplace_us_0_update_0_stage_69;
  reg [31:0] dark_laplace_us_0_update_0_stage_70;
  reg [31:0] dark_laplace_us_0_update_0_stage_71;
  reg [31:0] dark_laplace_us_0_update_0_stage_72;
  reg [31:0] dark_laplace_us_0_update_0_stage_73;
  reg [31:0] dark_laplace_us_0_update_0_stage_74;
  reg [31:0] dark_laplace_us_0_update_0_stage_75;
  reg [31:0] dark_laplace_us_0_update_0_stage_76;
  reg [31:0] dark_laplace_us_0_update_0_stage_77;
  reg [31:0] dark_laplace_us_0_update_0_stage_78;
  reg [31:0] dark_laplace_us_0_update_0_stage_79;
  reg [31:0] dark_laplace_us_0_update_0_stage_80;
  reg [31:0] dark_laplace_us_0_update_0_stage_81;
  reg [31:0] dark_laplace_us_0_update_0_stage_82;
  reg [31:0] dark_laplace_us_0_update_0_stage_83;
  reg [31:0] dark_laplace_us_0_update_0_stage_84;
  reg [31:0] dark_laplace_us_0_update_0_stage_85;
  reg [31:0] dark_laplace_us_0_update_0_stage_86;
  reg [31:0] dark_laplace_us_0_update_0_stage_87;
  reg [31:0] dark_laplace_us_0_update_0_stage_88;
  reg [31:0] dark_laplace_us_0_update_0_stage_89;
  reg [31:0] dark_laplace_us_0_update_0_stage_90;
  reg [31:0] dark_laplace_us_0_update_0_stage_91;
  reg [31:0] dark_laplace_us_0_update_0_stage_92;
  reg [31:0] dark_laplace_us_0_update_0_stage_93;
  reg [31:0] dark_laplace_us_0_update_0_stage_94;
  reg [31:0] dark_laplace_us_0_update_0_stage_95;
  reg [31:0] dark_laplace_us_0_update_0_stage_96;
  reg [31:0] dark_laplace_us_0_update_0_stage_97;
  reg [31:0] dark_laplace_us_0_update_0_stage_98;
  reg [31:0] dark_laplace_us_0_update_0_stage_99;
  reg [31:0] dark_laplace_us_0_update_0_stage_100;
  reg [31:0] dark_laplace_us_0_update_0_stage_101;
  reg [31:0] dark_laplace_us_0_update_0_stage_102;
  reg [31:0] dark_laplace_us_0_update_0_stage_103;
  reg [31:0] dark_laplace_us_0_update_0_stage_104;
  reg [31:0] dark_laplace_us_0_update_0_stage_105;
  reg [31:0] dark_laplace_us_0_update_0_stage_106;
  reg [31:0] dark_laplace_us_0_update_0_stage_107;
  reg [31:0] dark_laplace_us_0_update_0_stage_108;
  reg [31:0] dark_laplace_us_0_update_0_stage_109;
  reg [31:0] dark_laplace_us_0_update_0_stage_110;
  reg [31:0] dark_laplace_us_0_update_0_stage_111;
  reg [31:0] dark_laplace_us_0_update_0_stage_112;
  reg [31:0] dark_laplace_us_0_update_0_stage_113;
  reg [31:0] dark_laplace_us_0_update_0_stage_114;
  reg [31:0] dark_laplace_us_0_update_0_stage_115;
  reg [31:0] dark_laplace_us_0_update_0_stage_116;
  reg [31:0] dark_laplace_us_0_update_0_stage_117;
  reg [31:0] dark_laplace_us_0_update_0_stage_118;
  reg [31:0] dark_laplace_us_0_update_0_stage_119;
  reg [31:0] dark_laplace_us_0_update_0_stage_120;
  reg [31:0] dark_laplace_us_0_update_0_stage_121;
  reg [31:0] dark_laplace_us_0_update_0_stage_122;
  reg [31:0] dark_laplace_us_0_update_0_stage_123;
  reg [31:0] dark_laplace_us_0_update_0_stage_124;
  reg [31:0] dark_laplace_us_0_update_0_stage_125;
  reg [31:0] dark_laplace_us_0_update_0_stage_126;
  reg [31:0] dark_laplace_us_0_update_0_stage_127;
  reg [31:0] dark_laplace_us_0_update_0_stage_128;
  reg [31:0] dark_laplace_us_0_update_0_stage_129;
  reg [31:0] dark_laplace_us_0_update_0_stage_130;
  reg [31:0] dark_laplace_us_0_update_0_stage_131;
  reg [31:0] dark_laplace_us_0_update_0_stage_132;
  reg [31:0] dark_laplace_us_0_update_0_stage_133;
  reg [31:0] dark_laplace_us_0_update_0_stage_134;
  reg [31:0] dark_laplace_us_0_update_0_stage_135;
  reg [31:0] dark_laplace_us_0_update_0_stage_136;
  reg [31:0] dark_laplace_us_0_update_0_stage_137;
  reg [31:0] dark_laplace_us_0_update_0_stage_138;
  reg [31:0] dark_laplace_us_0_update_0_stage_139;
  reg [31:0] dark_laplace_us_0_update_0_stage_140;
  reg [31:0] dark_laplace_us_0_update_0_stage_141;
  reg [31:0] dark_laplace_us_0_update_0_stage_142;
  reg [31:0] dark_laplace_us_0_update_0_stage_143;
  reg [31:0] dark_laplace_us_0_update_0_stage_144;
  reg [31:0] dark_laplace_us_0_update_0_stage_145;
  reg [31:0] dark_laplace_us_0_update_0_stage_146;
  reg [31:0] dark_laplace_us_0_update_0_stage_147;
  reg [31:0] dark_laplace_us_0_update_0_stage_148;
  reg [31:0] dark_laplace_us_0_update_0_stage_149;
  reg [31:0] dark_laplace_us_0_update_0_stage_150;
  reg [31:0] dark_laplace_us_0_update_0_stage_151;
  reg [31:0] dark_laplace_us_0_update_0_stage_152;
  reg [31:0] dark_laplace_us_0_update_0_stage_153;
  reg [31:0] dark_laplace_us_0_update_0_stage_154;
  reg [31:0] dark_laplace_us_0_update_0_stage_155;
  reg [31:0] dark_laplace_us_0_update_0_stage_156;
  reg [31:0] dark_laplace_us_0_update_0_stage_157;
  reg [31:0] dark_laplace_us_0_update_0_stage_158;
  reg [31:0] dark_laplace_us_0_update_0_stage_159;
  reg [31:0] dark_laplace_us_0_update_0_stage_160;
  reg [31:0] dark_laplace_us_0_update_0_stage_161;
  reg [31:0] dark_laplace_us_0_update_0_stage_162;
  reg [31:0] dark_laplace_us_0_update_0_stage_163;
  reg [31:0] dark_laplace_us_0_update_0_stage_164;
  reg [31:0] dark_laplace_us_0_update_0_stage_165;
  reg [31:0] dark_laplace_us_0_update_0_stage_166;
  reg [31:0] dark_laplace_us_0_update_0_stage_167;
  reg [31:0] dark_laplace_us_0_update_0_stage_168;
  reg [31:0] dark_laplace_us_0_update_0_stage_169;
  reg [31:0] dark_laplace_us_0_update_0_stage_170;
  reg [31:0] dark_laplace_us_0_update_0_stage_171;
  reg [31:0] dark_laplace_us_0_update_0_stage_172;
  reg [31:0] dark_laplace_us_0_update_0_stage_173;
  reg [31:0] dark_laplace_us_0_update_0_stage_174;
  reg [31:0] dark_laplace_us_0_update_0_stage_175;
  reg [31:0] dark_laplace_us_0_update_0_stage_176;
  reg [31:0] dark_laplace_us_0_update_0_stage_177;
  reg [31:0] dark_laplace_us_0_update_0_stage_178;
  reg [31:0] dark_laplace_us_0_update_0_stage_179;
  reg [31:0] dark_laplace_us_0_update_0_stage_180;
  reg [31:0] dark_laplace_us_0_update_0_stage_181;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_28;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_29;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_30;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_31;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_32;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_33;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_34;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_35;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_36;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_37;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_38;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_39;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_40;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_41;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_42;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_43;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_44;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_45;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_46;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_47;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_48;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_49;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_50;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_51;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_52;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_53;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_54;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_55;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_56;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_57;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_58;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_59;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_60;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_61;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_62;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_63;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_64;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_65;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_66;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_67;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_68;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_69;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_70;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_71;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_72;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_73;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_74;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_75;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_76;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_77;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_78;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_79;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_80;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_81;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_82;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_83;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_84;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_85;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_86;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_87;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_88;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_89;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_90;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_91;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_92;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_93;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_94;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_95;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_96;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_97;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_98;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_99;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_100;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_101;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_102;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_103;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_104;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_105;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_106;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_107;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_108;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_109;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_110;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_111;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_112;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_113;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_114;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_115;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_116;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_117;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_118;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_119;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_120;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_121;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_122;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_123;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_124;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_125;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_126;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_127;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_128;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_129;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_130;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_131;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_132;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_133;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_134;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_135;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_136;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_137;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_138;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_139;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_140;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_141;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_142;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_143;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_144;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_145;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_146;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_147;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_148;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_149;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_150;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_151;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_152;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_153;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_154;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_155;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_156;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_157;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_158;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_159;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_160;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_161;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_162;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_163;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_164;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_165;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_166;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_167;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_168;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_169;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_170;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_171;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_172;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_173;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_174;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_175;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_176;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_177;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_178;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_179;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_180;
  reg [31:0] dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_181;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_35;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_36;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_37;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_38;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_39;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_40;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_41;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_42;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_43;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_44;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_45;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_46;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_47;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_48;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_49;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_50;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_51;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_52;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_53;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_54;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_55;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_56;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_57;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_58;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_59;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_60;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_61;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_62;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_63;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_64;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_65;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_66;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_67;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_68;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_69;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_70;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_71;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_72;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_73;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_74;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_75;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_76;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_77;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_78;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_79;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_80;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_81;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_82;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_83;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_84;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_85;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_86;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_87;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_88;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_89;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_90;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_91;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_92;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_93;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_94;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_95;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_96;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_97;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_98;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_99;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_100;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_101;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_102;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_103;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_104;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_105;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_106;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_107;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_108;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_109;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_110;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_111;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_112;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_113;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_114;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_115;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_116;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_117;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_118;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_119;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_120;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_121;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_122;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_123;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_124;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_125;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_126;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_127;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_128;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_129;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_130;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_131;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_132;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_133;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_134;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_135;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_136;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_137;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_138;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_139;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_140;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_141;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_142;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_143;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_144;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_145;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_146;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_147;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_148;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_149;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_150;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_151;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_152;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_153;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_154;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_155;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_156;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_157;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_158;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_159;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_160;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_161;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_162;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_163;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_164;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_165;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_166;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_167;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_168;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_169;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_170;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_171;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_172;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_173;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_174;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_175;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_176;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_177;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_178;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_179;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_180;
  reg [31:0] dark_weights_weight_sums_update_0_read_read_22_stage_181;
  reg [31:0] weight_sums_update_0_stage_37;
  reg [31:0] weight_sums_update_0_stage_38;
  reg [31:0] weight_sums_update_0_stage_39;
  reg [31:0] weight_sums_update_0_stage_40;
  reg [31:0] weight_sums_update_0_stage_41;
  reg [31:0] weight_sums_update_0_stage_42;
  reg [31:0] weight_sums_update_0_stage_43;
  reg [31:0] weight_sums_update_0_stage_44;
  reg [31:0] weight_sums_update_0_stage_45;
  reg [31:0] weight_sums_update_0_stage_46;
  reg [31:0] weight_sums_update_0_stage_47;
  reg [31:0] weight_sums_update_0_stage_48;
  reg [31:0] weight_sums_update_0_stage_49;
  reg [31:0] weight_sums_update_0_stage_50;
  reg [31:0] weight_sums_update_0_stage_51;
  reg [31:0] weight_sums_update_0_stage_52;
  reg [31:0] weight_sums_update_0_stage_53;
  reg [31:0] weight_sums_update_0_stage_54;
  reg [31:0] weight_sums_update_0_stage_55;
  reg [31:0] weight_sums_update_0_stage_56;
  reg [31:0] weight_sums_update_0_stage_57;
  reg [31:0] weight_sums_update_0_stage_58;
  reg [31:0] weight_sums_update_0_stage_59;
  reg [31:0] weight_sums_update_0_stage_60;
  reg [31:0] weight_sums_update_0_stage_61;
  reg [31:0] weight_sums_update_0_stage_62;
  reg [31:0] weight_sums_update_0_stage_63;
  reg [31:0] weight_sums_update_0_stage_64;
  reg [31:0] weight_sums_update_0_stage_65;
  reg [31:0] weight_sums_update_0_stage_66;
  reg [31:0] weight_sums_update_0_stage_67;
  reg [31:0] weight_sums_update_0_stage_68;
  reg [31:0] weight_sums_update_0_stage_69;
  reg [31:0] weight_sums_update_0_stage_70;
  reg [31:0] weight_sums_update_0_stage_71;
  reg [31:0] weight_sums_update_0_stage_72;
  reg [31:0] weight_sums_update_0_stage_73;
  reg [31:0] weight_sums_update_0_stage_74;
  reg [31:0] weight_sums_update_0_stage_75;
  reg [31:0] weight_sums_update_0_stage_76;
  reg [31:0] weight_sums_update_0_stage_77;
  reg [31:0] weight_sums_update_0_stage_78;
  reg [31:0] weight_sums_update_0_stage_79;
  reg [31:0] weight_sums_update_0_stage_80;
  reg [31:0] weight_sums_update_0_stage_81;
  reg [31:0] weight_sums_update_0_stage_82;
  reg [31:0] weight_sums_update_0_stage_83;
  reg [31:0] weight_sums_update_0_stage_84;
  reg [31:0] weight_sums_update_0_stage_85;
  reg [31:0] weight_sums_update_0_stage_86;
  reg [31:0] weight_sums_update_0_stage_87;
  reg [31:0] weight_sums_update_0_stage_88;
  reg [31:0] weight_sums_update_0_stage_89;
  reg [31:0] weight_sums_update_0_stage_90;
  reg [31:0] weight_sums_update_0_stage_91;
  reg [31:0] weight_sums_update_0_stage_92;
  reg [31:0] weight_sums_update_0_stage_93;
  reg [31:0] weight_sums_update_0_stage_94;
  reg [31:0] weight_sums_update_0_stage_95;
  reg [31:0] weight_sums_update_0_stage_96;
  reg [31:0] weight_sums_update_0_stage_97;
  reg [31:0] weight_sums_update_0_stage_98;
  reg [31:0] weight_sums_update_0_stage_99;
  reg [31:0] weight_sums_update_0_stage_100;
  reg [31:0] weight_sums_update_0_stage_101;
  reg [31:0] weight_sums_update_0_stage_102;
  reg [31:0] weight_sums_update_0_stage_103;
  reg [31:0] weight_sums_update_0_stage_104;
  reg [31:0] weight_sums_update_0_stage_105;
  reg [31:0] weight_sums_update_0_stage_106;
  reg [31:0] weight_sums_update_0_stage_107;
  reg [31:0] weight_sums_update_0_stage_108;
  reg [31:0] weight_sums_update_0_stage_109;
  reg [31:0] weight_sums_update_0_stage_110;
  reg [31:0] weight_sums_update_0_stage_111;
  reg [31:0] weight_sums_update_0_stage_112;
  reg [31:0] weight_sums_update_0_stage_113;
  reg [31:0] weight_sums_update_0_stage_114;
  reg [31:0] weight_sums_update_0_stage_115;
  reg [31:0] weight_sums_update_0_stage_116;
  reg [31:0] weight_sums_update_0_stage_117;
  reg [31:0] weight_sums_update_0_stage_118;
  reg [31:0] weight_sums_update_0_stage_119;
  reg [31:0] weight_sums_update_0_stage_120;
  reg [31:0] weight_sums_update_0_stage_121;
  reg [31:0] weight_sums_update_0_stage_122;
  reg [31:0] weight_sums_update_0_stage_123;
  reg [31:0] weight_sums_update_0_stage_124;
  reg [31:0] weight_sums_update_0_stage_125;
  reg [31:0] weight_sums_update_0_stage_126;
  reg [31:0] weight_sums_update_0_stage_127;
  reg [31:0] weight_sums_update_0_stage_128;
  reg [31:0] weight_sums_update_0_stage_129;
  reg [31:0] weight_sums_update_0_stage_130;
  reg [31:0] weight_sums_update_0_stage_131;
  reg [31:0] weight_sums_update_0_stage_132;
  reg [31:0] weight_sums_update_0_stage_133;
  reg [31:0] weight_sums_update_0_stage_134;
  reg [31:0] weight_sums_update_0_stage_135;
  reg [31:0] weight_sums_update_0_stage_136;
  reg [31:0] weight_sums_update_0_stage_137;
  reg [31:0] weight_sums_update_0_stage_138;
  reg [31:0] weight_sums_update_0_stage_139;
  reg [31:0] weight_sums_update_0_stage_140;
  reg [31:0] weight_sums_update_0_stage_141;
  reg [31:0] weight_sums_update_0_stage_142;
  reg [31:0] weight_sums_update_0_stage_143;
  reg [31:0] weight_sums_update_0_stage_144;
  reg [31:0] weight_sums_update_0_stage_145;
  reg [31:0] weight_sums_update_0_stage_146;
  reg [31:0] weight_sums_update_0_stage_147;
  reg [31:0] weight_sums_update_0_stage_148;
  reg [31:0] weight_sums_update_0_stage_149;
  reg [31:0] weight_sums_update_0_stage_150;
  reg [31:0] weight_sums_update_0_stage_151;
  reg [31:0] weight_sums_update_0_stage_152;
  reg [31:0] weight_sums_update_0_stage_153;
  reg [31:0] weight_sums_update_0_stage_154;
  reg [31:0] weight_sums_update_0_stage_155;
  reg [31:0] weight_sums_update_0_stage_156;
  reg [31:0] weight_sums_update_0_stage_157;
  reg [31:0] weight_sums_update_0_stage_158;
  reg [31:0] weight_sums_update_0_stage_159;
  reg [31:0] weight_sums_update_0_stage_160;
  reg [31:0] weight_sums_update_0_stage_161;
  reg [31:0] weight_sums_update_0_stage_162;
  reg [31:0] weight_sums_update_0_stage_163;
  reg [31:0] weight_sums_update_0_stage_164;
  reg [31:0] weight_sums_update_0_stage_165;
  reg [31:0] weight_sums_update_0_stage_166;
  reg [31:0] weight_sums_update_0_stage_167;
  reg [31:0] weight_sums_update_0_stage_168;
  reg [31:0] weight_sums_update_0_stage_169;
  reg [31:0] weight_sums_update_0_stage_170;
  reg [31:0] weight_sums_update_0_stage_171;
  reg [31:0] weight_sums_update_0_stage_172;
  reg [31:0] weight_sums_update_0_stage_173;
  reg [31:0] weight_sums_update_0_stage_174;
  reg [31:0] weight_sums_update_0_stage_175;
  reg [31:0] weight_sums_update_0_stage_176;
  reg [31:0] weight_sums_update_0_stage_177;
  reg [31:0] weight_sums_update_0_stage_178;
  reg [31:0] weight_sums_update_0_stage_179;
  reg [31:0] weight_sums_update_0_stage_180;
  reg [31:0] weight_sums_update_0_stage_181;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_36;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_37;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_38;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_39;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_40;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_41;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_42;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_43;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_44;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_45;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_46;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_47;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_48;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_49;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_50;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_51;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_52;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_53;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_54;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_55;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_56;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_57;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_58;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_59;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_60;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_61;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_62;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_63;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_64;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_65;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_66;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_67;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_68;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_69;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_70;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_71;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_72;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_73;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_74;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_75;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_76;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_77;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_78;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_79;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_80;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_81;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_82;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_83;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_84;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_85;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_86;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_87;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_88;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_89;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_90;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_91;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_92;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_93;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_94;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_95;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_96;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_97;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_98;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_99;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_100;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_101;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_102;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_103;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_104;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_105;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_106;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_107;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_108;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_109;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_110;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_111;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_112;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_113;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_114;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_115;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_116;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_117;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_118;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_119;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_120;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_121;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_122;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_123;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_124;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_125;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_126;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_127;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_128;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_129;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_130;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_131;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_132;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_133;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_134;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_135;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_136;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_137;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_138;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_139;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_140;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_141;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_142;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_143;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_144;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_145;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_146;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_147;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_148;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_149;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_150;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_151;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_152;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_153;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_154;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_155;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_156;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_157;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_158;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_159;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_160;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_161;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_162;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_163;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_164;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_165;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_166;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_167;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_168;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_169;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_170;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_171;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_172;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_173;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_174;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_175;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_176;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_177;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_178;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_179;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_180;
  reg [31:0] bright_weights_weight_sums_update_0_read_read_23_stage_181;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_38;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_39;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_40;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_41;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_42;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_43;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_44;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_45;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_46;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_47;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_48;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_49;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_50;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_51;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_52;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_53;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_54;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_55;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_56;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_57;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_58;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_59;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_60;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_61;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_62;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_63;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_64;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_65;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_66;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_67;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_68;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_69;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_70;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_71;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_72;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_73;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_74;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_75;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_76;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_77;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_78;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_79;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_80;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_81;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_82;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_83;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_84;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_85;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_86;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_87;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_88;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_89;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_90;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_91;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_92;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_93;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_94;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_95;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_96;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_97;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_98;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_99;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_100;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_101;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_102;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_103;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_104;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_105;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_106;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_107;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_108;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_109;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_110;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_111;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_112;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_113;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_114;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_115;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_116;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_117;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_118;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_119;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_120;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_121;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_122;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_123;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_124;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_125;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_126;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_127;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_128;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_129;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_130;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_131;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_132;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_133;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_134;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_135;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_136;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_137;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_138;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_139;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_140;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_141;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_142;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_143;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_144;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_145;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_146;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_147;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_148;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_149;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_150;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_151;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_152;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_153;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_154;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_155;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_156;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_157;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_158;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_159;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_160;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_161;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_162;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_163;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_164;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_165;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_166;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_167;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_168;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_169;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_170;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_171;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_172;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_173;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_174;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_175;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_176;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_177;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_178;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_179;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_180;
  reg [31:0] weight_sums_weight_sums_update_0_write_write_24_stage_181;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_42;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_43;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_44;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_45;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_46;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_47;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_48;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_49;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_50;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_51;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_52;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_53;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_54;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_55;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_56;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_57;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_58;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_59;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_60;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_61;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_62;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_63;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_64;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_65;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_66;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_67;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_68;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_69;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_70;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_71;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_72;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_73;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_74;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_75;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_76;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_77;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_78;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_79;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_80;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_81;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_82;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_83;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_84;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_85;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_86;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_87;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_88;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_89;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_90;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_91;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_92;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_93;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_94;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_95;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_96;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_97;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_98;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_99;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_100;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_101;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_102;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_103;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_104;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_105;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_106;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_107;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_108;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_109;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_110;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_111;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_112;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_113;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_114;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_115;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_116;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_117;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_118;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_119;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_120;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_121;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_122;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_123;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_124;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_125;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_126;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_127;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_128;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_129;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_130;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_131;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_132;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_133;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_134;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_135;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_136;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_137;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_138;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_139;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_140;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_141;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_142;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_143;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_144;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_145;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_146;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_147;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_148;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_149;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_150;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_151;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_152;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_153;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_154;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_155;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_156;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_157;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_158;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_159;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_160;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_161;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_162;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_163;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_164;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_165;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_166;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_167;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_168;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_169;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_170;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_171;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_172;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_173;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_174;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_175;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_176;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_177;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_178;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_179;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_180;
  reg [31:0] dark_dark_laplace_diff_0_update_0_read_read_27_stage_181;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_43;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_44;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_45;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_46;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_47;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_48;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_49;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_50;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_51;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_52;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_53;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_54;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_55;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_56;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_57;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_58;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_59;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_60;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_61;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_62;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_63;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_64;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_65;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_66;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_67;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_68;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_69;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_70;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_71;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_72;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_73;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_74;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_75;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_76;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_77;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_78;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_79;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_80;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_81;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_82;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_83;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_84;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_85;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_86;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_87;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_88;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_89;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_90;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_91;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_92;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_93;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_94;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_95;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_96;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_97;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_98;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_99;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_100;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_101;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_102;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_103;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_104;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_105;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_106;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_107;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_108;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_109;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_110;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_111;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_112;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_113;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_114;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_115;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_116;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_117;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_118;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_119;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_120;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_121;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_122;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_123;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_124;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_125;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_126;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_127;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_128;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_129;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_130;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_131;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_132;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_133;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_134;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_135;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_136;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_137;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_138;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_139;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_140;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_141;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_142;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_143;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_144;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_145;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_146;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_147;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_148;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_149;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_150;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_151;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_152;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_153;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_154;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_155;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_156;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_157;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_158;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_159;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_160;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_161;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_162;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_163;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_164;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_165;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_166;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_167;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_168;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_169;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_170;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_171;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_172;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_173;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_174;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_175;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_176;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_177;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_178;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_179;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_180;
  reg [31:0] dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_181;
  reg [31:0] dark_laplace_diff_0_update_0_stage_44;
  reg [31:0] dark_laplace_diff_0_update_0_stage_45;
  reg [31:0] dark_laplace_diff_0_update_0_stage_46;
  reg [31:0] dark_laplace_diff_0_update_0_stage_47;
  reg [31:0] dark_laplace_diff_0_update_0_stage_48;
  reg [31:0] dark_laplace_diff_0_update_0_stage_49;
  reg [31:0] dark_laplace_diff_0_update_0_stage_50;
  reg [31:0] dark_laplace_diff_0_update_0_stage_51;
  reg [31:0] dark_laplace_diff_0_update_0_stage_52;
  reg [31:0] dark_laplace_diff_0_update_0_stage_53;
  reg [31:0] dark_laplace_diff_0_update_0_stage_54;
  reg [31:0] dark_laplace_diff_0_update_0_stage_55;
  reg [31:0] dark_laplace_diff_0_update_0_stage_56;
  reg [31:0] dark_laplace_diff_0_update_0_stage_57;
  reg [31:0] dark_laplace_diff_0_update_0_stage_58;
  reg [31:0] dark_laplace_diff_0_update_0_stage_59;
  reg [31:0] dark_laplace_diff_0_update_0_stage_60;
  reg [31:0] dark_laplace_diff_0_update_0_stage_61;
  reg [31:0] dark_laplace_diff_0_update_0_stage_62;
  reg [31:0] dark_laplace_diff_0_update_0_stage_63;
  reg [31:0] dark_laplace_diff_0_update_0_stage_64;
  reg [31:0] dark_laplace_diff_0_update_0_stage_65;
  reg [31:0] dark_laplace_diff_0_update_0_stage_66;
  reg [31:0] dark_laplace_diff_0_update_0_stage_67;
  reg [31:0] dark_laplace_diff_0_update_0_stage_68;
  reg [31:0] dark_laplace_diff_0_update_0_stage_69;
  reg [31:0] dark_laplace_diff_0_update_0_stage_70;
  reg [31:0] dark_laplace_diff_0_update_0_stage_71;
  reg [31:0] dark_laplace_diff_0_update_0_stage_72;
  reg [31:0] dark_laplace_diff_0_update_0_stage_73;
  reg [31:0] dark_laplace_diff_0_update_0_stage_74;
  reg [31:0] dark_laplace_diff_0_update_0_stage_75;
  reg [31:0] dark_laplace_diff_0_update_0_stage_76;
  reg [31:0] dark_laplace_diff_0_update_0_stage_77;
  reg [31:0] dark_laplace_diff_0_update_0_stage_78;
  reg [31:0] dark_laplace_diff_0_update_0_stage_79;
  reg [31:0] dark_laplace_diff_0_update_0_stage_80;
  reg [31:0] dark_laplace_diff_0_update_0_stage_81;
  reg [31:0] dark_laplace_diff_0_update_0_stage_82;
  reg [31:0] dark_laplace_diff_0_update_0_stage_83;
  reg [31:0] dark_laplace_diff_0_update_0_stage_84;
  reg [31:0] dark_laplace_diff_0_update_0_stage_85;
  reg [31:0] dark_laplace_diff_0_update_0_stage_86;
  reg [31:0] dark_laplace_diff_0_update_0_stage_87;
  reg [31:0] dark_laplace_diff_0_update_0_stage_88;
  reg [31:0] dark_laplace_diff_0_update_0_stage_89;
  reg [31:0] dark_laplace_diff_0_update_0_stage_90;
  reg [31:0] dark_laplace_diff_0_update_0_stage_91;
  reg [31:0] dark_laplace_diff_0_update_0_stage_92;
  reg [31:0] dark_laplace_diff_0_update_0_stage_93;
  reg [31:0] dark_laplace_diff_0_update_0_stage_94;
  reg [31:0] dark_laplace_diff_0_update_0_stage_95;
  reg [31:0] dark_laplace_diff_0_update_0_stage_96;
  reg [31:0] dark_laplace_diff_0_update_0_stage_97;
  reg [31:0] dark_laplace_diff_0_update_0_stage_98;
  reg [31:0] dark_laplace_diff_0_update_0_stage_99;
  reg [31:0] dark_laplace_diff_0_update_0_stage_100;
  reg [31:0] dark_laplace_diff_0_update_0_stage_101;
  reg [31:0] dark_laplace_diff_0_update_0_stage_102;
  reg [31:0] dark_laplace_diff_0_update_0_stage_103;
  reg [31:0] dark_laplace_diff_0_update_0_stage_104;
  reg [31:0] dark_laplace_diff_0_update_0_stage_105;
  reg [31:0] dark_laplace_diff_0_update_0_stage_106;
  reg [31:0] dark_laplace_diff_0_update_0_stage_107;
  reg [31:0] dark_laplace_diff_0_update_0_stage_108;
  reg [31:0] dark_laplace_diff_0_update_0_stage_109;
  reg [31:0] dark_laplace_diff_0_update_0_stage_110;
  reg [31:0] dark_laplace_diff_0_update_0_stage_111;
  reg [31:0] dark_laplace_diff_0_update_0_stage_112;
  reg [31:0] dark_laplace_diff_0_update_0_stage_113;
  reg [31:0] dark_laplace_diff_0_update_0_stage_114;
  reg [31:0] dark_laplace_diff_0_update_0_stage_115;
  reg [31:0] dark_laplace_diff_0_update_0_stage_116;
  reg [31:0] dark_laplace_diff_0_update_0_stage_117;
  reg [31:0] dark_laplace_diff_0_update_0_stage_118;
  reg [31:0] dark_laplace_diff_0_update_0_stage_119;
  reg [31:0] dark_laplace_diff_0_update_0_stage_120;
  reg [31:0] dark_laplace_diff_0_update_0_stage_121;
  reg [31:0] dark_laplace_diff_0_update_0_stage_122;
  reg [31:0] dark_laplace_diff_0_update_0_stage_123;
  reg [31:0] dark_laplace_diff_0_update_0_stage_124;
  reg [31:0] dark_laplace_diff_0_update_0_stage_125;
  reg [31:0] dark_laplace_diff_0_update_0_stage_126;
  reg [31:0] dark_laplace_diff_0_update_0_stage_127;
  reg [31:0] dark_laplace_diff_0_update_0_stage_128;
  reg [31:0] dark_laplace_diff_0_update_0_stage_129;
  reg [31:0] dark_laplace_diff_0_update_0_stage_130;
  reg [31:0] dark_laplace_diff_0_update_0_stage_131;
  reg [31:0] dark_laplace_diff_0_update_0_stage_132;
  reg [31:0] dark_laplace_diff_0_update_0_stage_133;
  reg [31:0] dark_laplace_diff_0_update_0_stage_134;
  reg [31:0] dark_laplace_diff_0_update_0_stage_135;
  reg [31:0] dark_laplace_diff_0_update_0_stage_136;
  reg [31:0] dark_laplace_diff_0_update_0_stage_137;
  reg [31:0] dark_laplace_diff_0_update_0_stage_138;
  reg [31:0] dark_laplace_diff_0_update_0_stage_139;
  reg [31:0] dark_laplace_diff_0_update_0_stage_140;
  reg [31:0] dark_laplace_diff_0_update_0_stage_141;
  reg [31:0] dark_laplace_diff_0_update_0_stage_142;
  reg [31:0] dark_laplace_diff_0_update_0_stage_143;
  reg [31:0] dark_laplace_diff_0_update_0_stage_144;
  reg [31:0] dark_laplace_diff_0_update_0_stage_145;
  reg [31:0] dark_laplace_diff_0_update_0_stage_146;
  reg [31:0] dark_laplace_diff_0_update_0_stage_147;
  reg [31:0] dark_laplace_diff_0_update_0_stage_148;
  reg [31:0] dark_laplace_diff_0_update_0_stage_149;
  reg [31:0] dark_laplace_diff_0_update_0_stage_150;
  reg [31:0] dark_laplace_diff_0_update_0_stage_151;
  reg [31:0] dark_laplace_diff_0_update_0_stage_152;
  reg [31:0] dark_laplace_diff_0_update_0_stage_153;
  reg [31:0] dark_laplace_diff_0_update_0_stage_154;
  reg [31:0] dark_laplace_diff_0_update_0_stage_155;
  reg [31:0] dark_laplace_diff_0_update_0_stage_156;
  reg [31:0] dark_laplace_diff_0_update_0_stage_157;
  reg [31:0] dark_laplace_diff_0_update_0_stage_158;
  reg [31:0] dark_laplace_diff_0_update_0_stage_159;
  reg [31:0] dark_laplace_diff_0_update_0_stage_160;
  reg [31:0] dark_laplace_diff_0_update_0_stage_161;
  reg [31:0] dark_laplace_diff_0_update_0_stage_162;
  reg [31:0] dark_laplace_diff_0_update_0_stage_163;
  reg [31:0] dark_laplace_diff_0_update_0_stage_164;
  reg [31:0] dark_laplace_diff_0_update_0_stage_165;
  reg [31:0] dark_laplace_diff_0_update_0_stage_166;
  reg [31:0] dark_laplace_diff_0_update_0_stage_167;
  reg [31:0] dark_laplace_diff_0_update_0_stage_168;
  reg [31:0] dark_laplace_diff_0_update_0_stage_169;
  reg [31:0] dark_laplace_diff_0_update_0_stage_170;
  reg [31:0] dark_laplace_diff_0_update_0_stage_171;
  reg [31:0] dark_laplace_diff_0_update_0_stage_172;
  reg [31:0] dark_laplace_diff_0_update_0_stage_173;
  reg [31:0] dark_laplace_diff_0_update_0_stage_174;
  reg [31:0] dark_laplace_diff_0_update_0_stage_175;
  reg [31:0] dark_laplace_diff_0_update_0_stage_176;
  reg [31:0] dark_laplace_diff_0_update_0_stage_177;
  reg [31:0] dark_laplace_diff_0_update_0_stage_178;
  reg [31:0] dark_laplace_diff_0_update_0_stage_179;
  reg [31:0] dark_laplace_diff_0_update_0_stage_180;
  reg [31:0] dark_laplace_diff_0_update_0_stage_181;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_45;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_46;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_47;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_48;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_49;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_50;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_51;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_52;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_53;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_54;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_55;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_56;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_57;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_58;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_59;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_60;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_61;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_62;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_63;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_64;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_65;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_66;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_67;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_68;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_69;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_70;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_71;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_72;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_73;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_74;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_75;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_76;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_77;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_78;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_79;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_80;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_81;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_82;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_83;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_84;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_85;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_86;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_87;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_88;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_89;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_90;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_91;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_92;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_93;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_94;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_95;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_96;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_97;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_98;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_99;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_100;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_101;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_102;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_103;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_104;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_105;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_106;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_107;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_108;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_109;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_110;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_111;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_112;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_113;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_114;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_115;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_116;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_117;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_118;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_119;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_120;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_121;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_122;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_123;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_124;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_125;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_126;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_127;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_128;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_129;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_130;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_131;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_132;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_133;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_134;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_135;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_136;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_137;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_138;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_139;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_140;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_141;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_142;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_143;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_144;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_145;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_146;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_147;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_148;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_149;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_150;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_151;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_152;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_153;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_154;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_155;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_156;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_157;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_158;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_159;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_160;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_161;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_162;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_163;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_164;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_165;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_166;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_167;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_168;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_169;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_170;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_171;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_172;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_173;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_174;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_175;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_176;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_177;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_178;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_179;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_180;
  reg [31:0] dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_181;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_49;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_50;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_51;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_52;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_53;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_54;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_55;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_56;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_57;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_58;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_59;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_60;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_61;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_62;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_63;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_64;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_65;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_66;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_67;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_68;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_69;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_70;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_71;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_72;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_73;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_74;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_75;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_76;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_77;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_78;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_79;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_80;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_81;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_82;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_83;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_84;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_85;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_86;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_87;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_88;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_89;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_90;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_91;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_92;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_93;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_94;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_95;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_96;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_97;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_98;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_99;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_100;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_101;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_102;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_103;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_104;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_105;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_106;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_107;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_108;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_109;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_110;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_111;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_112;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_113;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_114;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_115;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_116;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_117;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_118;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_119;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_120;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_121;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_122;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_123;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_124;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_125;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_126;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_127;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_128;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_129;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_130;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_131;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_132;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_133;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_134;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_135;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_136;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_137;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_138;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_139;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_140;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_141;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_142;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_143;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_144;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_145;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_146;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_147;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_148;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_149;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_150;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_151;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_152;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_153;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_154;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_155;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_156;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_157;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_158;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_159;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_160;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_161;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_162;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_163;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_164;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_165;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_166;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_167;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_168;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_169;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_170;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_171;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_172;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_173;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_174;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_175;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_176;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_177;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_178;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_179;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_180;
  reg [31:0] bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_181;
  reg [31:0] bright_gauss_ds_2_update_0_stage_50;
  reg [31:0] bright_gauss_ds_2_update_0_stage_51;
  reg [31:0] bright_gauss_ds_2_update_0_stage_52;
  reg [31:0] bright_gauss_ds_2_update_0_stage_53;
  reg [31:0] bright_gauss_ds_2_update_0_stage_54;
  reg [31:0] bright_gauss_ds_2_update_0_stage_55;
  reg [31:0] bright_gauss_ds_2_update_0_stage_56;
  reg [31:0] bright_gauss_ds_2_update_0_stage_57;
  reg [31:0] bright_gauss_ds_2_update_0_stage_58;
  reg [31:0] bright_gauss_ds_2_update_0_stage_59;
  reg [31:0] bright_gauss_ds_2_update_0_stage_60;
  reg [31:0] bright_gauss_ds_2_update_0_stage_61;
  reg [31:0] bright_gauss_ds_2_update_0_stage_62;
  reg [31:0] bright_gauss_ds_2_update_0_stage_63;
  reg [31:0] bright_gauss_ds_2_update_0_stage_64;
  reg [31:0] bright_gauss_ds_2_update_0_stage_65;
  reg [31:0] bright_gauss_ds_2_update_0_stage_66;
  reg [31:0] bright_gauss_ds_2_update_0_stage_67;
  reg [31:0] bright_gauss_ds_2_update_0_stage_68;
  reg [31:0] bright_gauss_ds_2_update_0_stage_69;
  reg [31:0] bright_gauss_ds_2_update_0_stage_70;
  reg [31:0] bright_gauss_ds_2_update_0_stage_71;
  reg [31:0] bright_gauss_ds_2_update_0_stage_72;
  reg [31:0] bright_gauss_ds_2_update_0_stage_73;
  reg [31:0] bright_gauss_ds_2_update_0_stage_74;
  reg [31:0] bright_gauss_ds_2_update_0_stage_75;
  reg [31:0] bright_gauss_ds_2_update_0_stage_76;
  reg [31:0] bright_gauss_ds_2_update_0_stage_77;
  reg [31:0] bright_gauss_ds_2_update_0_stage_78;
  reg [31:0] bright_gauss_ds_2_update_0_stage_79;
  reg [31:0] bright_gauss_ds_2_update_0_stage_80;
  reg [31:0] bright_gauss_ds_2_update_0_stage_81;
  reg [31:0] bright_gauss_ds_2_update_0_stage_82;
  reg [31:0] bright_gauss_ds_2_update_0_stage_83;
  reg [31:0] bright_gauss_ds_2_update_0_stage_84;
  reg [31:0] bright_gauss_ds_2_update_0_stage_85;
  reg [31:0] bright_gauss_ds_2_update_0_stage_86;
  reg [31:0] bright_gauss_ds_2_update_0_stage_87;
  reg [31:0] bright_gauss_ds_2_update_0_stage_88;
  reg [31:0] bright_gauss_ds_2_update_0_stage_89;
  reg [31:0] bright_gauss_ds_2_update_0_stage_90;
  reg [31:0] bright_gauss_ds_2_update_0_stage_91;
  reg [31:0] bright_gauss_ds_2_update_0_stage_92;
  reg [31:0] bright_gauss_ds_2_update_0_stage_93;
  reg [31:0] bright_gauss_ds_2_update_0_stage_94;
  reg [31:0] bright_gauss_ds_2_update_0_stage_95;
  reg [31:0] bright_gauss_ds_2_update_0_stage_96;
  reg [31:0] bright_gauss_ds_2_update_0_stage_97;
  reg [31:0] bright_gauss_ds_2_update_0_stage_98;
  reg [31:0] bright_gauss_ds_2_update_0_stage_99;
  reg [31:0] bright_gauss_ds_2_update_0_stage_100;
  reg [31:0] bright_gauss_ds_2_update_0_stage_101;
  reg [31:0] bright_gauss_ds_2_update_0_stage_102;
  reg [31:0] bright_gauss_ds_2_update_0_stage_103;
  reg [31:0] bright_gauss_ds_2_update_0_stage_104;
  reg [31:0] bright_gauss_ds_2_update_0_stage_105;
  reg [31:0] bright_gauss_ds_2_update_0_stage_106;
  reg [31:0] bright_gauss_ds_2_update_0_stage_107;
  reg [31:0] bright_gauss_ds_2_update_0_stage_108;
  reg [31:0] bright_gauss_ds_2_update_0_stage_109;
  reg [31:0] bright_gauss_ds_2_update_0_stage_110;
  reg [31:0] bright_gauss_ds_2_update_0_stage_111;
  reg [31:0] bright_gauss_ds_2_update_0_stage_112;
  reg [31:0] bright_gauss_ds_2_update_0_stage_113;
  reg [31:0] bright_gauss_ds_2_update_0_stage_114;
  reg [31:0] bright_gauss_ds_2_update_0_stage_115;
  reg [31:0] bright_gauss_ds_2_update_0_stage_116;
  reg [31:0] bright_gauss_ds_2_update_0_stage_117;
  reg [31:0] bright_gauss_ds_2_update_0_stage_118;
  reg [31:0] bright_gauss_ds_2_update_0_stage_119;
  reg [31:0] bright_gauss_ds_2_update_0_stage_120;
  reg [31:0] bright_gauss_ds_2_update_0_stage_121;
  reg [31:0] bright_gauss_ds_2_update_0_stage_122;
  reg [31:0] bright_gauss_ds_2_update_0_stage_123;
  reg [31:0] bright_gauss_ds_2_update_0_stage_124;
  reg [31:0] bright_gauss_ds_2_update_0_stage_125;
  reg [31:0] bright_gauss_ds_2_update_0_stage_126;
  reg [31:0] bright_gauss_ds_2_update_0_stage_127;
  reg [31:0] bright_gauss_ds_2_update_0_stage_128;
  reg [31:0] bright_gauss_ds_2_update_0_stage_129;
  reg [31:0] bright_gauss_ds_2_update_0_stage_130;
  reg [31:0] bright_gauss_ds_2_update_0_stage_131;
  reg [31:0] bright_gauss_ds_2_update_0_stage_132;
  reg [31:0] bright_gauss_ds_2_update_0_stage_133;
  reg [31:0] bright_gauss_ds_2_update_0_stage_134;
  reg [31:0] bright_gauss_ds_2_update_0_stage_135;
  reg [31:0] bright_gauss_ds_2_update_0_stage_136;
  reg [31:0] bright_gauss_ds_2_update_0_stage_137;
  reg [31:0] bright_gauss_ds_2_update_0_stage_138;
  reg [31:0] bright_gauss_ds_2_update_0_stage_139;
  reg [31:0] bright_gauss_ds_2_update_0_stage_140;
  reg [31:0] bright_gauss_ds_2_update_0_stage_141;
  reg [31:0] bright_gauss_ds_2_update_0_stage_142;
  reg [31:0] bright_gauss_ds_2_update_0_stage_143;
  reg [31:0] bright_gauss_ds_2_update_0_stage_144;
  reg [31:0] bright_gauss_ds_2_update_0_stage_145;
  reg [31:0] bright_gauss_ds_2_update_0_stage_146;
  reg [31:0] bright_gauss_ds_2_update_0_stage_147;
  reg [31:0] bright_gauss_ds_2_update_0_stage_148;
  reg [31:0] bright_gauss_ds_2_update_0_stage_149;
  reg [31:0] bright_gauss_ds_2_update_0_stage_150;
  reg [31:0] bright_gauss_ds_2_update_0_stage_151;
  reg [31:0] bright_gauss_ds_2_update_0_stage_152;
  reg [31:0] bright_gauss_ds_2_update_0_stage_153;
  reg [31:0] bright_gauss_ds_2_update_0_stage_154;
  reg [31:0] bright_gauss_ds_2_update_0_stage_155;
  reg [31:0] bright_gauss_ds_2_update_0_stage_156;
  reg [31:0] bright_gauss_ds_2_update_0_stage_157;
  reg [31:0] bright_gauss_ds_2_update_0_stage_158;
  reg [31:0] bright_gauss_ds_2_update_0_stage_159;
  reg [31:0] bright_gauss_ds_2_update_0_stage_160;
  reg [31:0] bright_gauss_ds_2_update_0_stage_161;
  reg [31:0] bright_gauss_ds_2_update_0_stage_162;
  reg [31:0] bright_gauss_ds_2_update_0_stage_163;
  reg [31:0] bright_gauss_ds_2_update_0_stage_164;
  reg [31:0] bright_gauss_ds_2_update_0_stage_165;
  reg [31:0] bright_gauss_ds_2_update_0_stage_166;
  reg [31:0] bright_gauss_ds_2_update_0_stage_167;
  reg [31:0] bright_gauss_ds_2_update_0_stage_168;
  reg [31:0] bright_gauss_ds_2_update_0_stage_169;
  reg [31:0] bright_gauss_ds_2_update_0_stage_170;
  reg [31:0] bright_gauss_ds_2_update_0_stage_171;
  reg [31:0] bright_gauss_ds_2_update_0_stage_172;
  reg [31:0] bright_gauss_ds_2_update_0_stage_173;
  reg [31:0] bright_gauss_ds_2_update_0_stage_174;
  reg [31:0] bright_gauss_ds_2_update_0_stage_175;
  reg [31:0] bright_gauss_ds_2_update_0_stage_176;
  reg [31:0] bright_gauss_ds_2_update_0_stage_177;
  reg [31:0] bright_gauss_ds_2_update_0_stage_178;
  reg [31:0] bright_gauss_ds_2_update_0_stage_179;
  reg [31:0] bright_gauss_ds_2_update_0_stage_180;
  reg [31:0] bright_gauss_ds_2_update_0_stage_181;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_58;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_59;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_60;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_61;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_62;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_63;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_64;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_65;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_66;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_67;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_68;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_69;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_70;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_71;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_72;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_73;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_74;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_75;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_76;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_77;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_78;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_79;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_80;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_81;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_82;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_83;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_84;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_85;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_86;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_87;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_88;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_89;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_90;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_91;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_92;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_93;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_94;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_95;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_96;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_97;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_98;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_99;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_100;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_101;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_102;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_103;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_104;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_105;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_106;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_107;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_108;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_109;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_110;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_111;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_112;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_113;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_114;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_115;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_116;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_117;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_118;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_119;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_120;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_121;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_122;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_123;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_124;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_125;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_126;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_127;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_128;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_129;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_130;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_131;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_132;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_133;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_134;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_135;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_136;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_137;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_138;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_139;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_140;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_141;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_142;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_143;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_144;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_145;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_146;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_147;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_148;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_149;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_150;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_151;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_152;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_153;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_154;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_155;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_156;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_157;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_158;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_159;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_160;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_161;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_162;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_163;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_164;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_165;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_166;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_167;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_168;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_169;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_170;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_171;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_172;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_173;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_174;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_175;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_176;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_177;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_178;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_179;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_180;
  reg [31:0] bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_181;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_51;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_52;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_53;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_54;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_55;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_56;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_57;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_58;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_59;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_60;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_61;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_62;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_63;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_64;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_65;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_66;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_67;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_68;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_69;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_70;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_71;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_72;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_73;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_74;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_75;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_76;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_77;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_78;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_79;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_80;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_81;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_82;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_83;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_84;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_85;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_86;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_87;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_88;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_89;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_90;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_91;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_92;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_93;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_94;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_95;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_96;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_97;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_98;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_99;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_100;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_101;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_102;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_103;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_104;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_105;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_106;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_107;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_108;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_109;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_110;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_111;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_112;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_113;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_114;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_115;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_116;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_117;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_118;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_119;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_120;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_121;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_122;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_123;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_124;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_125;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_126;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_127;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_128;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_129;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_130;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_131;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_132;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_133;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_134;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_135;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_136;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_137;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_138;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_139;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_140;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_141;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_142;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_143;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_144;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_145;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_146;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_147;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_148;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_149;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_150;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_151;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_152;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_153;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_154;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_155;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_156;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_157;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_158;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_159;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_160;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_161;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_162;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_163;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_164;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_165;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_166;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_167;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_168;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_169;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_170;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_171;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_172;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_173;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_174;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_175;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_176;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_177;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_178;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_179;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_180;
  reg [31:0] bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_181;
  reg [31:0] bright_gauss_ds_3_update_0_stage_59;
  reg [31:0] bright_gauss_ds_3_update_0_stage_60;
  reg [31:0] bright_gauss_ds_3_update_0_stage_61;
  reg [31:0] bright_gauss_ds_3_update_0_stage_62;
  reg [31:0] bright_gauss_ds_3_update_0_stage_63;
  reg [31:0] bright_gauss_ds_3_update_0_stage_64;
  reg [31:0] bright_gauss_ds_3_update_0_stage_65;
  reg [31:0] bright_gauss_ds_3_update_0_stage_66;
  reg [31:0] bright_gauss_ds_3_update_0_stage_67;
  reg [31:0] bright_gauss_ds_3_update_0_stage_68;
  reg [31:0] bright_gauss_ds_3_update_0_stage_69;
  reg [31:0] bright_gauss_ds_3_update_0_stage_70;
  reg [31:0] bright_gauss_ds_3_update_0_stage_71;
  reg [31:0] bright_gauss_ds_3_update_0_stage_72;
  reg [31:0] bright_gauss_ds_3_update_0_stage_73;
  reg [31:0] bright_gauss_ds_3_update_0_stage_74;
  reg [31:0] bright_gauss_ds_3_update_0_stage_75;
  reg [31:0] bright_gauss_ds_3_update_0_stage_76;
  reg [31:0] bright_gauss_ds_3_update_0_stage_77;
  reg [31:0] bright_gauss_ds_3_update_0_stage_78;
  reg [31:0] bright_gauss_ds_3_update_0_stage_79;
  reg [31:0] bright_gauss_ds_3_update_0_stage_80;
  reg [31:0] bright_gauss_ds_3_update_0_stage_81;
  reg [31:0] bright_gauss_ds_3_update_0_stage_82;
  reg [31:0] bright_gauss_ds_3_update_0_stage_83;
  reg [31:0] bright_gauss_ds_3_update_0_stage_84;
  reg [31:0] bright_gauss_ds_3_update_0_stage_85;
  reg [31:0] bright_gauss_ds_3_update_0_stage_86;
  reg [31:0] bright_gauss_ds_3_update_0_stage_87;
  reg [31:0] bright_gauss_ds_3_update_0_stage_88;
  reg [31:0] bright_gauss_ds_3_update_0_stage_89;
  reg [31:0] bright_gauss_ds_3_update_0_stage_90;
  reg [31:0] bright_gauss_ds_3_update_0_stage_91;
  reg [31:0] bright_gauss_ds_3_update_0_stage_92;
  reg [31:0] bright_gauss_ds_3_update_0_stage_93;
  reg [31:0] bright_gauss_ds_3_update_0_stage_94;
  reg [31:0] bright_gauss_ds_3_update_0_stage_95;
  reg [31:0] bright_gauss_ds_3_update_0_stage_96;
  reg [31:0] bright_gauss_ds_3_update_0_stage_97;
  reg [31:0] bright_gauss_ds_3_update_0_stage_98;
  reg [31:0] bright_gauss_ds_3_update_0_stage_99;
  reg [31:0] bright_gauss_ds_3_update_0_stage_100;
  reg [31:0] bright_gauss_ds_3_update_0_stage_101;
  reg [31:0] bright_gauss_ds_3_update_0_stage_102;
  reg [31:0] bright_gauss_ds_3_update_0_stage_103;
  reg [31:0] bright_gauss_ds_3_update_0_stage_104;
  reg [31:0] bright_gauss_ds_3_update_0_stage_105;
  reg [31:0] bright_gauss_ds_3_update_0_stage_106;
  reg [31:0] bright_gauss_ds_3_update_0_stage_107;
  reg [31:0] bright_gauss_ds_3_update_0_stage_108;
  reg [31:0] bright_gauss_ds_3_update_0_stage_109;
  reg [31:0] bright_gauss_ds_3_update_0_stage_110;
  reg [31:0] bright_gauss_ds_3_update_0_stage_111;
  reg [31:0] bright_gauss_ds_3_update_0_stage_112;
  reg [31:0] bright_gauss_ds_3_update_0_stage_113;
  reg [31:0] bright_gauss_ds_3_update_0_stage_114;
  reg [31:0] bright_gauss_ds_3_update_0_stage_115;
  reg [31:0] bright_gauss_ds_3_update_0_stage_116;
  reg [31:0] bright_gauss_ds_3_update_0_stage_117;
  reg [31:0] bright_gauss_ds_3_update_0_stage_118;
  reg [31:0] bright_gauss_ds_3_update_0_stage_119;
  reg [31:0] bright_gauss_ds_3_update_0_stage_120;
  reg [31:0] bright_gauss_ds_3_update_0_stage_121;
  reg [31:0] bright_gauss_ds_3_update_0_stage_122;
  reg [31:0] bright_gauss_ds_3_update_0_stage_123;
  reg [31:0] bright_gauss_ds_3_update_0_stage_124;
  reg [31:0] bright_gauss_ds_3_update_0_stage_125;
  reg [31:0] bright_gauss_ds_3_update_0_stage_126;
  reg [31:0] bright_gauss_ds_3_update_0_stage_127;
  reg [31:0] bright_gauss_ds_3_update_0_stage_128;
  reg [31:0] bright_gauss_ds_3_update_0_stage_129;
  reg [31:0] bright_gauss_ds_3_update_0_stage_130;
  reg [31:0] bright_gauss_ds_3_update_0_stage_131;
  reg [31:0] bright_gauss_ds_3_update_0_stage_132;
  reg [31:0] bright_gauss_ds_3_update_0_stage_133;
  reg [31:0] bright_gauss_ds_3_update_0_stage_134;
  reg [31:0] bright_gauss_ds_3_update_0_stage_135;
  reg [31:0] bright_gauss_ds_3_update_0_stage_136;
  reg [31:0] bright_gauss_ds_3_update_0_stage_137;
  reg [31:0] bright_gauss_ds_3_update_0_stage_138;
  reg [31:0] bright_gauss_ds_3_update_0_stage_139;
  reg [31:0] bright_gauss_ds_3_update_0_stage_140;
  reg [31:0] bright_gauss_ds_3_update_0_stage_141;
  reg [31:0] bright_gauss_ds_3_update_0_stage_142;
  reg [31:0] bright_gauss_ds_3_update_0_stage_143;
  reg [31:0] bright_gauss_ds_3_update_0_stage_144;
  reg [31:0] bright_gauss_ds_3_update_0_stage_145;
  reg [31:0] bright_gauss_ds_3_update_0_stage_146;
  reg [31:0] bright_gauss_ds_3_update_0_stage_147;
  reg [31:0] bright_gauss_ds_3_update_0_stage_148;
  reg [31:0] bright_gauss_ds_3_update_0_stage_149;
  reg [31:0] bright_gauss_ds_3_update_0_stage_150;
  reg [31:0] bright_gauss_ds_3_update_0_stage_151;
  reg [31:0] bright_gauss_ds_3_update_0_stage_152;
  reg [31:0] bright_gauss_ds_3_update_0_stage_153;
  reg [31:0] bright_gauss_ds_3_update_0_stage_154;
  reg [31:0] bright_gauss_ds_3_update_0_stage_155;
  reg [31:0] bright_gauss_ds_3_update_0_stage_156;
  reg [31:0] bright_gauss_ds_3_update_0_stage_157;
  reg [31:0] bright_gauss_ds_3_update_0_stage_158;
  reg [31:0] bright_gauss_ds_3_update_0_stage_159;
  reg [31:0] bright_gauss_ds_3_update_0_stage_160;
  reg [31:0] bright_gauss_ds_3_update_0_stage_161;
  reg [31:0] bright_gauss_ds_3_update_0_stage_162;
  reg [31:0] bright_gauss_ds_3_update_0_stage_163;
  reg [31:0] bright_gauss_ds_3_update_0_stage_164;
  reg [31:0] bright_gauss_ds_3_update_0_stage_165;
  reg [31:0] bright_gauss_ds_3_update_0_stage_166;
  reg [31:0] bright_gauss_ds_3_update_0_stage_167;
  reg [31:0] bright_gauss_ds_3_update_0_stage_168;
  reg [31:0] bright_gauss_ds_3_update_0_stage_169;
  reg [31:0] bright_gauss_ds_3_update_0_stage_170;
  reg [31:0] bright_gauss_ds_3_update_0_stage_171;
  reg [31:0] bright_gauss_ds_3_update_0_stage_172;
  reg [31:0] bright_gauss_ds_3_update_0_stage_173;
  reg [31:0] bright_gauss_ds_3_update_0_stage_174;
  reg [31:0] bright_gauss_ds_3_update_0_stage_175;
  reg [31:0] bright_gauss_ds_3_update_0_stage_176;
  reg [31:0] bright_gauss_ds_3_update_0_stage_177;
  reg [31:0] bright_gauss_ds_3_update_0_stage_178;
  reg [31:0] bright_gauss_ds_3_update_0_stage_179;
  reg [31:0] bright_gauss_ds_3_update_0_stage_180;
  reg [31:0] bright_gauss_ds_3_update_0_stage_181;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_64;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_65;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_66;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_67;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_68;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_69;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_70;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_71;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_72;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_73;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_74;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_75;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_76;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_77;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_78;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_79;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_80;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_81;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_82;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_83;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_84;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_85;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_86;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_87;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_88;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_89;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_90;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_91;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_92;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_93;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_94;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_95;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_96;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_97;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_98;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_99;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_100;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_101;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_102;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_103;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_104;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_105;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_106;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_107;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_108;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_109;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_110;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_111;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_112;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_113;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_114;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_115;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_116;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_117;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_118;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_119;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_120;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_121;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_122;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_123;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_124;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_125;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_126;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_127;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_128;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_129;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_130;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_131;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_132;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_133;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_134;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_135;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_136;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_137;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_138;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_139;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_140;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_141;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_142;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_143;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_144;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_145;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_146;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_147;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_148;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_149;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_150;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_151;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_152;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_153;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_154;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_155;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_156;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_157;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_158;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_159;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_160;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_161;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_162;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_163;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_164;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_165;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_166;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_167;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_168;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_169;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_170;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_171;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_172;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_173;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_174;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_175;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_176;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_177;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_178;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_179;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_180;
  reg [31:0] bright_bright_laplace_diff_0_update_0_read_read_42_stage_181;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_65;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_66;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_67;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_68;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_69;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_70;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_71;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_72;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_73;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_74;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_75;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_76;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_77;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_78;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_79;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_80;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_81;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_82;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_83;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_84;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_85;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_86;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_87;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_88;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_89;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_90;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_91;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_92;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_93;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_94;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_95;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_96;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_97;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_98;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_99;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_100;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_101;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_102;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_103;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_104;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_105;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_106;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_107;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_108;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_109;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_110;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_111;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_112;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_113;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_114;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_115;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_116;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_117;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_118;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_119;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_120;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_121;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_122;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_123;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_124;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_125;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_126;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_127;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_128;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_129;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_130;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_131;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_132;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_133;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_134;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_135;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_136;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_137;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_138;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_139;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_140;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_141;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_142;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_143;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_144;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_145;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_146;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_147;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_148;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_149;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_150;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_151;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_152;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_153;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_154;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_155;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_156;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_157;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_158;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_159;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_160;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_161;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_162;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_163;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_164;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_165;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_166;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_167;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_168;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_169;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_170;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_171;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_172;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_173;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_174;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_175;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_176;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_177;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_178;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_179;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_180;
  reg [31:0] bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_181;
  reg [31:0] bright_laplace_diff_0_update_0_stage_66;
  reg [31:0] bright_laplace_diff_0_update_0_stage_67;
  reg [31:0] bright_laplace_diff_0_update_0_stage_68;
  reg [31:0] bright_laplace_diff_0_update_0_stage_69;
  reg [31:0] bright_laplace_diff_0_update_0_stage_70;
  reg [31:0] bright_laplace_diff_0_update_0_stage_71;
  reg [31:0] bright_laplace_diff_0_update_0_stage_72;
  reg [31:0] bright_laplace_diff_0_update_0_stage_73;
  reg [31:0] bright_laplace_diff_0_update_0_stage_74;
  reg [31:0] bright_laplace_diff_0_update_0_stage_75;
  reg [31:0] bright_laplace_diff_0_update_0_stage_76;
  reg [31:0] bright_laplace_diff_0_update_0_stage_77;
  reg [31:0] bright_laplace_diff_0_update_0_stage_78;
  reg [31:0] bright_laplace_diff_0_update_0_stage_79;
  reg [31:0] bright_laplace_diff_0_update_0_stage_80;
  reg [31:0] bright_laplace_diff_0_update_0_stage_81;
  reg [31:0] bright_laplace_diff_0_update_0_stage_82;
  reg [31:0] bright_laplace_diff_0_update_0_stage_83;
  reg [31:0] bright_laplace_diff_0_update_0_stage_84;
  reg [31:0] bright_laplace_diff_0_update_0_stage_85;
  reg [31:0] bright_laplace_diff_0_update_0_stage_86;
  reg [31:0] bright_laplace_diff_0_update_0_stage_87;
  reg [31:0] bright_laplace_diff_0_update_0_stage_88;
  reg [31:0] bright_laplace_diff_0_update_0_stage_89;
  reg [31:0] bright_laplace_diff_0_update_0_stage_90;
  reg [31:0] bright_laplace_diff_0_update_0_stage_91;
  reg [31:0] bright_laplace_diff_0_update_0_stage_92;
  reg [31:0] bright_laplace_diff_0_update_0_stage_93;
  reg [31:0] bright_laplace_diff_0_update_0_stage_94;
  reg [31:0] bright_laplace_diff_0_update_0_stage_95;
  reg [31:0] bright_laplace_diff_0_update_0_stage_96;
  reg [31:0] bright_laplace_diff_0_update_0_stage_97;
  reg [31:0] bright_laplace_diff_0_update_0_stage_98;
  reg [31:0] bright_laplace_diff_0_update_0_stage_99;
  reg [31:0] bright_laplace_diff_0_update_0_stage_100;
  reg [31:0] bright_laplace_diff_0_update_0_stage_101;
  reg [31:0] bright_laplace_diff_0_update_0_stage_102;
  reg [31:0] bright_laplace_diff_0_update_0_stage_103;
  reg [31:0] bright_laplace_diff_0_update_0_stage_104;
  reg [31:0] bright_laplace_diff_0_update_0_stage_105;
  reg [31:0] bright_laplace_diff_0_update_0_stage_106;
  reg [31:0] bright_laplace_diff_0_update_0_stage_107;
  reg [31:0] bright_laplace_diff_0_update_0_stage_108;
  reg [31:0] bright_laplace_diff_0_update_0_stage_109;
  reg [31:0] bright_laplace_diff_0_update_0_stage_110;
  reg [31:0] bright_laplace_diff_0_update_0_stage_111;
  reg [31:0] bright_laplace_diff_0_update_0_stage_112;
  reg [31:0] bright_laplace_diff_0_update_0_stage_113;
  reg [31:0] bright_laplace_diff_0_update_0_stage_114;
  reg [31:0] bright_laplace_diff_0_update_0_stage_115;
  reg [31:0] bright_laplace_diff_0_update_0_stage_116;
  reg [31:0] bright_laplace_diff_0_update_0_stage_117;
  reg [31:0] bright_laplace_diff_0_update_0_stage_118;
  reg [31:0] bright_laplace_diff_0_update_0_stage_119;
  reg [31:0] bright_laplace_diff_0_update_0_stage_120;
  reg [31:0] bright_laplace_diff_0_update_0_stage_121;
  reg [31:0] bright_laplace_diff_0_update_0_stage_122;
  reg [31:0] bright_laplace_diff_0_update_0_stage_123;
  reg [31:0] bright_laplace_diff_0_update_0_stage_124;
  reg [31:0] bright_laplace_diff_0_update_0_stage_125;
  reg [31:0] bright_laplace_diff_0_update_0_stage_126;
  reg [31:0] bright_laplace_diff_0_update_0_stage_127;
  reg [31:0] bright_laplace_diff_0_update_0_stage_128;
  reg [31:0] bright_laplace_diff_0_update_0_stage_129;
  reg [31:0] bright_laplace_diff_0_update_0_stage_130;
  reg [31:0] bright_laplace_diff_0_update_0_stage_131;
  reg [31:0] bright_laplace_diff_0_update_0_stage_132;
  reg [31:0] bright_laplace_diff_0_update_0_stage_133;
  reg [31:0] bright_laplace_diff_0_update_0_stage_134;
  reg [31:0] bright_laplace_diff_0_update_0_stage_135;
  reg [31:0] bright_laplace_diff_0_update_0_stage_136;
  reg [31:0] bright_laplace_diff_0_update_0_stage_137;
  reg [31:0] bright_laplace_diff_0_update_0_stage_138;
  reg [31:0] bright_laplace_diff_0_update_0_stage_139;
  reg [31:0] bright_laplace_diff_0_update_0_stage_140;
  reg [31:0] bright_laplace_diff_0_update_0_stage_141;
  reg [31:0] bright_laplace_diff_0_update_0_stage_142;
  reg [31:0] bright_laplace_diff_0_update_0_stage_143;
  reg [31:0] bright_laplace_diff_0_update_0_stage_144;
  reg [31:0] bright_laplace_diff_0_update_0_stage_145;
  reg [31:0] bright_laplace_diff_0_update_0_stage_146;
  reg [31:0] bright_laplace_diff_0_update_0_stage_147;
  reg [31:0] bright_laplace_diff_0_update_0_stage_148;
  reg [31:0] bright_laplace_diff_0_update_0_stage_149;
  reg [31:0] bright_laplace_diff_0_update_0_stage_150;
  reg [31:0] bright_laplace_diff_0_update_0_stage_151;
  reg [31:0] bright_laplace_diff_0_update_0_stage_152;
  reg [31:0] bright_laplace_diff_0_update_0_stage_153;
  reg [31:0] bright_laplace_diff_0_update_0_stage_154;
  reg [31:0] bright_laplace_diff_0_update_0_stage_155;
  reg [31:0] bright_laplace_diff_0_update_0_stage_156;
  reg [31:0] bright_laplace_diff_0_update_0_stage_157;
  reg [31:0] bright_laplace_diff_0_update_0_stage_158;
  reg [31:0] bright_laplace_diff_0_update_0_stage_159;
  reg [31:0] bright_laplace_diff_0_update_0_stage_160;
  reg [31:0] bright_laplace_diff_0_update_0_stage_161;
  reg [31:0] bright_laplace_diff_0_update_0_stage_162;
  reg [31:0] bright_laplace_diff_0_update_0_stage_163;
  reg [31:0] bright_laplace_diff_0_update_0_stage_164;
  reg [31:0] bright_laplace_diff_0_update_0_stage_165;
  reg [31:0] bright_laplace_diff_0_update_0_stage_166;
  reg [31:0] bright_laplace_diff_0_update_0_stage_167;
  reg [31:0] bright_laplace_diff_0_update_0_stage_168;
  reg [31:0] bright_laplace_diff_0_update_0_stage_169;
  reg [31:0] bright_laplace_diff_0_update_0_stage_170;
  reg [31:0] bright_laplace_diff_0_update_0_stage_171;
  reg [31:0] bright_laplace_diff_0_update_0_stage_172;
  reg [31:0] bright_laplace_diff_0_update_0_stage_173;
  reg [31:0] bright_laplace_diff_0_update_0_stage_174;
  reg [31:0] bright_laplace_diff_0_update_0_stage_175;
  reg [31:0] bright_laplace_diff_0_update_0_stage_176;
  reg [31:0] bright_laplace_diff_0_update_0_stage_177;
  reg [31:0] bright_laplace_diff_0_update_0_stage_178;
  reg [31:0] bright_laplace_diff_0_update_0_stage_179;
  reg [31:0] bright_laplace_diff_0_update_0_stage_180;
  reg [31:0] bright_laplace_diff_0_update_0_stage_181;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_67;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_68;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_69;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_70;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_71;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_72;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_73;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_74;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_75;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_76;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_77;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_78;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_79;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_80;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_81;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_82;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_83;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_84;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_85;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_86;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_87;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_88;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_89;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_90;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_91;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_92;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_93;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_94;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_95;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_96;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_97;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_98;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_99;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_100;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_101;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_102;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_103;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_104;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_105;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_106;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_107;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_108;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_109;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_110;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_111;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_112;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_113;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_114;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_115;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_116;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_117;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_118;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_119;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_120;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_121;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_122;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_123;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_124;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_125;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_126;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_127;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_128;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_129;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_130;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_131;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_132;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_133;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_134;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_135;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_136;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_137;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_138;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_139;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_140;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_141;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_142;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_143;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_144;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_145;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_146;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_147;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_148;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_149;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_150;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_151;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_152;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_153;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_154;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_155;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_156;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_157;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_158;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_159;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_160;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_161;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_162;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_163;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_164;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_165;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_166;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_167;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_168;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_169;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_170;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_171;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_172;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_173;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_174;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_175;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_176;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_177;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_178;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_179;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_180;
  reg [31:0] bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_181;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_72;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_73;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_74;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_75;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_76;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_77;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_78;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_79;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_80;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_81;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_82;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_83;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_84;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_85;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_86;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_87;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_88;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_89;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_90;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_91;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_92;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_93;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_94;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_95;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_96;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_97;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_98;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_99;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_100;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_101;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_102;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_103;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_104;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_105;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_106;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_107;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_108;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_109;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_110;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_111;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_112;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_113;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_114;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_115;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_116;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_117;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_118;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_119;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_120;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_121;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_122;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_123;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_124;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_125;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_126;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_127;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_128;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_129;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_130;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_131;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_132;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_133;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_134;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_135;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_136;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_137;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_138;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_139;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_140;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_141;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_142;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_143;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_144;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_145;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_146;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_147;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_148;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_149;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_150;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_151;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_152;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_153;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_154;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_155;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_156;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_157;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_158;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_159;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_160;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_161;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_162;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_163;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_164;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_165;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_166;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_167;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_168;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_169;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_170;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_171;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_172;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_173;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_174;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_175;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_176;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_177;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_178;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_179;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_180;
  reg [31:0] bright_weights_bright_weights_normed_update_0_read_read_48_stage_181;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_73;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_74;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_75;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_76;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_77;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_78;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_79;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_80;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_81;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_82;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_83;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_84;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_85;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_86;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_87;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_88;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_89;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_90;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_91;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_92;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_93;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_94;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_95;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_96;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_97;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_98;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_99;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_100;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_101;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_102;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_103;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_104;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_105;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_106;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_107;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_108;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_109;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_110;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_111;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_112;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_113;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_114;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_115;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_116;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_117;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_118;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_119;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_120;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_121;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_122;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_123;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_124;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_125;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_126;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_127;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_128;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_129;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_130;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_131;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_132;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_133;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_134;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_135;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_136;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_137;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_138;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_139;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_140;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_141;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_142;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_143;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_144;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_145;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_146;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_147;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_148;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_149;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_150;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_151;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_152;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_153;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_154;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_155;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_156;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_157;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_158;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_159;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_160;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_161;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_162;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_163;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_164;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_165;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_166;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_167;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_168;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_169;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_170;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_171;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_172;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_173;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_174;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_175;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_176;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_177;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_178;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_179;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_180;
  reg [31:0] weight_sums_bright_weights_normed_update_0_read_read_49_stage_181;
  reg [31:0] bright_weights_normed_update_0_stage_74;
  reg [31:0] bright_weights_normed_update_0_stage_75;
  reg [31:0] bright_weights_normed_update_0_stage_76;
  reg [31:0] bright_weights_normed_update_0_stage_77;
  reg [31:0] bright_weights_normed_update_0_stage_78;
  reg [31:0] bright_weights_normed_update_0_stage_79;
  reg [31:0] bright_weights_normed_update_0_stage_80;
  reg [31:0] bright_weights_normed_update_0_stage_81;
  reg [31:0] bright_weights_normed_update_0_stage_82;
  reg [31:0] bright_weights_normed_update_0_stage_83;
  reg [31:0] bright_weights_normed_update_0_stage_84;
  reg [31:0] bright_weights_normed_update_0_stage_85;
  reg [31:0] bright_weights_normed_update_0_stage_86;
  reg [31:0] bright_weights_normed_update_0_stage_87;
  reg [31:0] bright_weights_normed_update_0_stage_88;
  reg [31:0] bright_weights_normed_update_0_stage_89;
  reg [31:0] bright_weights_normed_update_0_stage_90;
  reg [31:0] bright_weights_normed_update_0_stage_91;
  reg [31:0] bright_weights_normed_update_0_stage_92;
  reg [31:0] bright_weights_normed_update_0_stage_93;
  reg [31:0] bright_weights_normed_update_0_stage_94;
  reg [31:0] bright_weights_normed_update_0_stage_95;
  reg [31:0] bright_weights_normed_update_0_stage_96;
  reg [31:0] bright_weights_normed_update_0_stage_97;
  reg [31:0] bright_weights_normed_update_0_stage_98;
  reg [31:0] bright_weights_normed_update_0_stage_99;
  reg [31:0] bright_weights_normed_update_0_stage_100;
  reg [31:0] bright_weights_normed_update_0_stage_101;
  reg [31:0] bright_weights_normed_update_0_stage_102;
  reg [31:0] bright_weights_normed_update_0_stage_103;
  reg [31:0] bright_weights_normed_update_0_stage_104;
  reg [31:0] bright_weights_normed_update_0_stage_105;
  reg [31:0] bright_weights_normed_update_0_stage_106;
  reg [31:0] bright_weights_normed_update_0_stage_107;
  reg [31:0] bright_weights_normed_update_0_stage_108;
  reg [31:0] bright_weights_normed_update_0_stage_109;
  reg [31:0] bright_weights_normed_update_0_stage_110;
  reg [31:0] bright_weights_normed_update_0_stage_111;
  reg [31:0] bright_weights_normed_update_0_stage_112;
  reg [31:0] bright_weights_normed_update_0_stage_113;
  reg [31:0] bright_weights_normed_update_0_stage_114;
  reg [31:0] bright_weights_normed_update_0_stage_115;
  reg [31:0] bright_weights_normed_update_0_stage_116;
  reg [31:0] bright_weights_normed_update_0_stage_117;
  reg [31:0] bright_weights_normed_update_0_stage_118;
  reg [31:0] bright_weights_normed_update_0_stage_119;
  reg [31:0] bright_weights_normed_update_0_stage_120;
  reg [31:0] bright_weights_normed_update_0_stage_121;
  reg [31:0] bright_weights_normed_update_0_stage_122;
  reg [31:0] bright_weights_normed_update_0_stage_123;
  reg [31:0] bright_weights_normed_update_0_stage_124;
  reg [31:0] bright_weights_normed_update_0_stage_125;
  reg [31:0] bright_weights_normed_update_0_stage_126;
  reg [31:0] bright_weights_normed_update_0_stage_127;
  reg [31:0] bright_weights_normed_update_0_stage_128;
  reg [31:0] bright_weights_normed_update_0_stage_129;
  reg [31:0] bright_weights_normed_update_0_stage_130;
  reg [31:0] bright_weights_normed_update_0_stage_131;
  reg [31:0] bright_weights_normed_update_0_stage_132;
  reg [31:0] bright_weights_normed_update_0_stage_133;
  reg [31:0] bright_weights_normed_update_0_stage_134;
  reg [31:0] bright_weights_normed_update_0_stage_135;
  reg [31:0] bright_weights_normed_update_0_stage_136;
  reg [31:0] bright_weights_normed_update_0_stage_137;
  reg [31:0] bright_weights_normed_update_0_stage_138;
  reg [31:0] bright_weights_normed_update_0_stage_139;
  reg [31:0] bright_weights_normed_update_0_stage_140;
  reg [31:0] bright_weights_normed_update_0_stage_141;
  reg [31:0] bright_weights_normed_update_0_stage_142;
  reg [31:0] bright_weights_normed_update_0_stage_143;
  reg [31:0] bright_weights_normed_update_0_stage_144;
  reg [31:0] bright_weights_normed_update_0_stage_145;
  reg [31:0] bright_weights_normed_update_0_stage_146;
  reg [31:0] bright_weights_normed_update_0_stage_147;
  reg [31:0] bright_weights_normed_update_0_stage_148;
  reg [31:0] bright_weights_normed_update_0_stage_149;
  reg [31:0] bright_weights_normed_update_0_stage_150;
  reg [31:0] bright_weights_normed_update_0_stage_151;
  reg [31:0] bright_weights_normed_update_0_stage_152;
  reg [31:0] bright_weights_normed_update_0_stage_153;
  reg [31:0] bright_weights_normed_update_0_stage_154;
  reg [31:0] bright_weights_normed_update_0_stage_155;
  reg [31:0] bright_weights_normed_update_0_stage_156;
  reg [31:0] bright_weights_normed_update_0_stage_157;
  reg [31:0] bright_weights_normed_update_0_stage_158;
  reg [31:0] bright_weights_normed_update_0_stage_159;
  reg [31:0] bright_weights_normed_update_0_stage_160;
  reg [31:0] bright_weights_normed_update_0_stage_161;
  reg [31:0] bright_weights_normed_update_0_stage_162;
  reg [31:0] bright_weights_normed_update_0_stage_163;
  reg [31:0] bright_weights_normed_update_0_stage_164;
  reg [31:0] bright_weights_normed_update_0_stage_165;
  reg [31:0] bright_weights_normed_update_0_stage_166;
  reg [31:0] bright_weights_normed_update_0_stage_167;
  reg [31:0] bright_weights_normed_update_0_stage_168;
  reg [31:0] bright_weights_normed_update_0_stage_169;
  reg [31:0] bright_weights_normed_update_0_stage_170;
  reg [31:0] bright_weights_normed_update_0_stage_171;
  reg [31:0] bright_weights_normed_update_0_stage_172;
  reg [31:0] bright_weights_normed_update_0_stage_173;
  reg [31:0] bright_weights_normed_update_0_stage_174;
  reg [31:0] bright_weights_normed_update_0_stage_175;
  reg [31:0] bright_weights_normed_update_0_stage_176;
  reg [31:0] bright_weights_normed_update_0_stage_177;
  reg [31:0] bright_weights_normed_update_0_stage_178;
  reg [31:0] bright_weights_normed_update_0_stage_179;
  reg [31:0] bright_weights_normed_update_0_stage_180;
  reg [31:0] bright_weights_normed_update_0_stage_181;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_75;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_76;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_77;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_78;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_79;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_80;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_81;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_82;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_83;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_84;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_85;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_86;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_87;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_88;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_89;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_90;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_91;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_92;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_93;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_94;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_95;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_96;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_97;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_98;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_99;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_100;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_101;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_102;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_103;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_104;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_105;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_106;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_107;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_108;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_109;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_110;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_111;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_112;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_113;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_114;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_115;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_116;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_117;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_118;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_119;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_120;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_121;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_122;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_123;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_124;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_125;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_126;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_127;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_128;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_129;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_130;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_131;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_132;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_133;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_134;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_135;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_136;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_137;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_138;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_139;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_140;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_141;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_142;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_143;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_144;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_145;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_146;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_147;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_148;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_149;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_150;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_151;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_152;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_153;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_154;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_155;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_156;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_157;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_158;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_159;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_160;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_161;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_162;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_163;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_164;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_165;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_166;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_167;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_168;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_169;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_170;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_171;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_172;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_173;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_174;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_175;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_176;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_177;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_178;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_179;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_180;
  reg [31:0] bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_79;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_80;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_81;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_82;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_83;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_84;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_85;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_86;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_87;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_88;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_89;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_90;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_91;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_92;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_93;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_80;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_81;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_82;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_83;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_84;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_85;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_86;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_87;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_88;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_89;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_90;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_91;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_92;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_93;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_94;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_95;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_96;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_97;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_98;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_99;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_100;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_101;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_102;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_103;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_104;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_105;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_106;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_107;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_108;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_109;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_110;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_111;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_112;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_113;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_114;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_115;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_116;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_117;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_118;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_119;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_120;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_121;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_122;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_123;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_124;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_125;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_126;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_127;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_128;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_129;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_130;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_131;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_132;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_133;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_134;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_135;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_136;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_1_update_0_stage_181;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_97;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_98;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_99;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_100;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_101;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_102;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_103;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_104;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_105;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_106;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_107;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_108;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_109;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_110;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_111;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_112;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_113;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_114;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_115;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_116;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_117;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_118;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_119;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_120;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_121;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_122;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_123;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_124;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_125;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_126;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_127;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_128;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_129;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_130;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_131;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_132;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_133;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_134;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_135;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_136;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_137;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_138;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_139;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_140;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_141;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_142;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_143;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_144;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_145;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_146;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_147;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_148;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_149;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_150;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_151;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_152;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_153;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_154;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_155;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_156;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_157;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_158;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_159;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_160;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_161;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_162;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_163;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_164;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_165;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_166;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_167;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_168;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_169;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_170;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_171;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_172;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_173;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_174;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_175;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_176;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_177;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_178;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_179;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_180;
  reg [287:0] dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_81;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_82;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_83;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_84;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_85;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_86;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_87;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_88;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_89;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_90;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_91;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_92;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_93;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_94;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_95;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_96;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_97;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_98;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_99;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_100;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_101;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_102;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_103;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_104;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_105;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_106;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_107;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_108;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_109;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_110;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_111;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_112;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_113;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_114;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_115;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_116;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_117;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_118;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_119;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_120;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_121;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_122;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_123;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_124;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_125;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_126;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_127;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_128;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_129;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_130;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_131;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_132;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_133;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_134;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_135;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_136;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_181;
  reg [31:0] dark_gauss_blur_3_update_0_stage_98;
  reg [31:0] dark_gauss_blur_3_update_0_stage_99;
  reg [31:0] dark_gauss_blur_3_update_0_stage_100;
  reg [31:0] dark_gauss_blur_3_update_0_stage_101;
  reg [31:0] dark_gauss_blur_3_update_0_stage_102;
  reg [31:0] dark_gauss_blur_3_update_0_stage_103;
  reg [31:0] dark_gauss_blur_3_update_0_stage_104;
  reg [31:0] dark_gauss_blur_3_update_0_stage_105;
  reg [31:0] dark_gauss_blur_3_update_0_stage_106;
  reg [31:0] dark_gauss_blur_3_update_0_stage_107;
  reg [31:0] dark_gauss_blur_3_update_0_stage_108;
  reg [31:0] dark_gauss_blur_3_update_0_stage_109;
  reg [31:0] dark_gauss_blur_3_update_0_stage_110;
  reg [31:0] dark_gauss_blur_3_update_0_stage_111;
  reg [31:0] dark_gauss_blur_3_update_0_stage_112;
  reg [31:0] dark_gauss_blur_3_update_0_stage_113;
  reg [31:0] dark_gauss_blur_3_update_0_stage_114;
  reg [31:0] dark_gauss_blur_3_update_0_stage_115;
  reg [31:0] dark_gauss_blur_3_update_0_stage_116;
  reg [31:0] dark_gauss_blur_3_update_0_stage_117;
  reg [31:0] dark_gauss_blur_3_update_0_stage_118;
  reg [31:0] dark_gauss_blur_3_update_0_stage_119;
  reg [31:0] dark_gauss_blur_3_update_0_stage_120;
  reg [31:0] dark_gauss_blur_3_update_0_stage_121;
  reg [31:0] dark_gauss_blur_3_update_0_stage_122;
  reg [31:0] dark_gauss_blur_3_update_0_stage_123;
  reg [31:0] dark_gauss_blur_3_update_0_stage_124;
  reg [31:0] dark_gauss_blur_3_update_0_stage_125;
  reg [31:0] dark_gauss_blur_3_update_0_stage_126;
  reg [31:0] dark_gauss_blur_3_update_0_stage_127;
  reg [31:0] dark_gauss_blur_3_update_0_stage_128;
  reg [31:0] dark_gauss_blur_3_update_0_stage_129;
  reg [31:0] dark_gauss_blur_3_update_0_stage_130;
  reg [31:0] dark_gauss_blur_3_update_0_stage_131;
  reg [31:0] dark_gauss_blur_3_update_0_stage_132;
  reg [31:0] dark_gauss_blur_3_update_0_stage_133;
  reg [31:0] dark_gauss_blur_3_update_0_stage_134;
  reg [31:0] dark_gauss_blur_3_update_0_stage_135;
  reg [31:0] dark_gauss_blur_3_update_0_stage_136;
  reg [31:0] dark_gauss_blur_3_update_0_stage_137;
  reg [31:0] dark_gauss_blur_3_update_0_stage_138;
  reg [31:0] dark_gauss_blur_3_update_0_stage_139;
  reg [31:0] dark_gauss_blur_3_update_0_stage_140;
  reg [31:0] dark_gauss_blur_3_update_0_stage_141;
  reg [31:0] dark_gauss_blur_3_update_0_stage_142;
  reg [31:0] dark_gauss_blur_3_update_0_stage_143;
  reg [31:0] dark_gauss_blur_3_update_0_stage_144;
  reg [31:0] dark_gauss_blur_3_update_0_stage_145;
  reg [31:0] dark_gauss_blur_3_update_0_stage_146;
  reg [31:0] dark_gauss_blur_3_update_0_stage_147;
  reg [31:0] dark_gauss_blur_3_update_0_stage_148;
  reg [31:0] dark_gauss_blur_3_update_0_stage_149;
  reg [31:0] dark_gauss_blur_3_update_0_stage_150;
  reg [31:0] dark_gauss_blur_3_update_0_stage_151;
  reg [31:0] dark_gauss_blur_3_update_0_stage_152;
  reg [31:0] dark_gauss_blur_3_update_0_stage_153;
  reg [31:0] dark_gauss_blur_3_update_0_stage_154;
  reg [31:0] dark_gauss_blur_3_update_0_stage_155;
  reg [31:0] dark_gauss_blur_3_update_0_stage_156;
  reg [31:0] dark_gauss_blur_3_update_0_stage_157;
  reg [31:0] dark_gauss_blur_3_update_0_stage_158;
  reg [31:0] dark_gauss_blur_3_update_0_stage_159;
  reg [31:0] dark_gauss_blur_3_update_0_stage_160;
  reg [31:0] dark_gauss_blur_3_update_0_stage_161;
  reg [31:0] dark_gauss_blur_3_update_0_stage_162;
  reg [31:0] dark_gauss_blur_3_update_0_stage_163;
  reg [31:0] dark_gauss_blur_3_update_0_stage_164;
  reg [31:0] dark_gauss_blur_3_update_0_stage_165;
  reg [31:0] dark_gauss_blur_3_update_0_stage_166;
  reg [31:0] dark_gauss_blur_3_update_0_stage_167;
  reg [31:0] dark_gauss_blur_3_update_0_stage_168;
  reg [31:0] dark_gauss_blur_3_update_0_stage_169;
  reg [31:0] dark_gauss_blur_3_update_0_stage_170;
  reg [31:0] dark_gauss_blur_3_update_0_stage_171;
  reg [31:0] dark_gauss_blur_3_update_0_stage_172;
  reg [31:0] dark_gauss_blur_3_update_0_stage_173;
  reg [31:0] dark_gauss_blur_3_update_0_stage_174;
  reg [31:0] dark_gauss_blur_3_update_0_stage_175;
  reg [31:0] dark_gauss_blur_3_update_0_stage_176;
  reg [31:0] dark_gauss_blur_3_update_0_stage_177;
  reg [31:0] dark_gauss_blur_3_update_0_stage_178;
  reg [31:0] dark_gauss_blur_3_update_0_stage_179;
  reg [31:0] dark_gauss_blur_3_update_0_stage_180;
  reg [31:0] dark_gauss_blur_3_update_0_stage_181;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_99;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_100;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_101;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_102;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_103;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_104;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_105;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_106;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_107;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_108;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_109;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_110;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_111;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_112;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_113;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_114;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_115;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_116;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_117;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_118;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_119;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_120;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_121;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_122;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_123;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_124;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_125;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_126;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_127;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_128;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_129;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_130;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_131;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_132;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_133;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_134;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_135;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_136;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_137;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_138;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_139;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_140;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_141;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_142;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_143;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_144;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_145;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_146;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_147;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_148;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_149;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_150;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_151;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_152;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_153;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_154;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_155;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_156;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_157;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_158;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_159;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_160;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_161;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_162;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_163;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_164;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_165;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_166;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_167;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_168;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_169;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_170;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_171;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_172;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_173;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_174;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_175;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_176;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_177;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_178;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_179;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_180;
  reg [31:0] dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_104;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_105;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_106;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_107;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_108;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_109;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_110;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_111;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_112;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_113;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_114;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_115;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_116;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_117;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_118;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_119;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_120;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_121;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_122;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_123;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_124;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_125;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_126;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_127;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_128;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_129;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_130;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_131;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_132;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_133;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_134;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_135;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_136;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_137;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_138;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_105;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_106;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_107;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_108;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_109;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_110;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_111;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_112;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_113;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_114;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_115;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_116;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_117;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_118;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_119;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_120;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_121;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_122;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_123;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_124;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_125;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_126;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_127;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_128;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_129;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_130;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_131;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_132;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_133;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_134;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_135;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_136;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_137;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_138;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_139;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_140;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_141;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_142;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_143;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_144;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_145;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_146;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_147;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_148;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_149;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_150;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_151;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_152;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_1_update_0_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_106;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_107;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_108;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_109;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_110;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_111;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_112;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_113;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_114;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_115;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_116;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_117;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_118;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_119;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_120;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_121;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_122;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_123;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_124;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_125;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_126;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_127;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_128;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_129;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_130;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_131;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_132;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_133;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_134;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_135;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_136;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_137;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_138;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_139;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_140;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_141;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_142;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_143;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_144;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_145;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_146;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_147;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_148;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_149;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_150;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_151;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_152;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_126;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_127;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_128;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_129;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_130;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_131;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_132;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_133;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_134;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_135;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_136;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_137;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_138;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_139;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_140;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_141;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_142;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_143;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_144;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_145;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_146;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_147;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_148;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_149;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_150;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_151;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_152;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_181;
  reg [31:0] fused_level_1_update_0_stage_128;
  reg [31:0] fused_level_1_update_0_stage_129;
  reg [31:0] fused_level_1_update_0_stage_130;
  reg [31:0] fused_level_1_update_0_stage_131;
  reg [31:0] fused_level_1_update_0_stage_132;
  reg [31:0] fused_level_1_update_0_stage_133;
  reg [31:0] fused_level_1_update_0_stage_134;
  reg [31:0] fused_level_1_update_0_stage_135;
  reg [31:0] fused_level_1_update_0_stage_136;
  reg [31:0] fused_level_1_update_0_stage_137;
  reg [31:0] fused_level_1_update_0_stage_138;
  reg [31:0] fused_level_1_update_0_stage_139;
  reg [31:0] fused_level_1_update_0_stage_140;
  reg [31:0] fused_level_1_update_0_stage_141;
  reg [31:0] fused_level_1_update_0_stage_142;
  reg [31:0] fused_level_1_update_0_stage_143;
  reg [31:0] fused_level_1_update_0_stage_144;
  reg [31:0] fused_level_1_update_0_stage_145;
  reg [31:0] fused_level_1_update_0_stage_146;
  reg [31:0] fused_level_1_update_0_stage_147;
  reg [31:0] fused_level_1_update_0_stage_148;
  reg [31:0] fused_level_1_update_0_stage_149;
  reg [31:0] fused_level_1_update_0_stage_150;
  reg [31:0] fused_level_1_update_0_stage_151;
  reg [31:0] fused_level_1_update_0_stage_152;
  reg [31:0] fused_level_1_update_0_stage_153;
  reg [31:0] fused_level_1_update_0_stage_154;
  reg [31:0] fused_level_1_update_0_stage_155;
  reg [31:0] fused_level_1_update_0_stage_156;
  reg [31:0] fused_level_1_update_0_stage_157;
  reg [31:0] fused_level_1_update_0_stage_158;
  reg [31:0] fused_level_1_update_0_stage_159;
  reg [31:0] fused_level_1_update_0_stage_160;
  reg [31:0] fused_level_1_update_0_stage_161;
  reg [31:0] fused_level_1_update_0_stage_162;
  reg [31:0] fused_level_1_update_0_stage_163;
  reg [31:0] fused_level_1_update_0_stage_164;
  reg [31:0] fused_level_1_update_0_stage_165;
  reg [31:0] fused_level_1_update_0_stage_166;
  reg [31:0] fused_level_1_update_0_stage_167;
  reg [31:0] fused_level_1_update_0_stage_168;
  reg [31:0] fused_level_1_update_0_stage_169;
  reg [31:0] fused_level_1_update_0_stage_170;
  reg [31:0] fused_level_1_update_0_stage_171;
  reg [31:0] fused_level_1_update_0_stage_172;
  reg [31:0] fused_level_1_update_0_stage_173;
  reg [31:0] fused_level_1_update_0_stage_174;
  reg [31:0] fused_level_1_update_0_stage_175;
  reg [31:0] fused_level_1_update_0_stage_176;
  reg [31:0] fused_level_1_update_0_stage_177;
  reg [31:0] fused_level_1_update_0_stage_178;
  reg [31:0] fused_level_1_update_0_stage_179;
  reg [31:0] fused_level_1_update_0_stage_180;
  reg [31:0] fused_level_1_update_0_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_127;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_128;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_129;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_130;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_131;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_132;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_133;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_134;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_135;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_136;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_181;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_129;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_130;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_131;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_132;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_133;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_134;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_135;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_136;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_137;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_138;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_139;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_140;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_141;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_142;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_143;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_144;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_145;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_146;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_147;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_148;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_149;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_150;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_151;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_152;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_153;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_154;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_155;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_156;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_157;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_158;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_159;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_160;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_161;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_162;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_163;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_164;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_165;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_166;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_167;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_168;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_169;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_170;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_171;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_172;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_173;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_174;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_175;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_176;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_177;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_178;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_179;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_180;
  reg [31:0] fused_level_1_fused_level_1_update_0_write_write_89_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_3_update_0_stage_181;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_142;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_143;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_144;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_145;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_146;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_147;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_148;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_149;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_150;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_151;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_152;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_153;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_154;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_155;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_156;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_157;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_158;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_159;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_160;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_161;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_162;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_163;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_164;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_165;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_166;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_167;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_168;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_169;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_170;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_171;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_172;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_173;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_174;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_175;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_176;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_177;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_178;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_179;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_180;
  reg [31:0] dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_181;
  reg [31:0] dark_laplace_us_2_update_0_stage_143;
  reg [31:0] dark_laplace_us_2_update_0_stage_144;
  reg [31:0] dark_laplace_us_2_update_0_stage_145;
  reg [31:0] dark_laplace_us_2_update_0_stage_146;
  reg [31:0] dark_laplace_us_2_update_0_stage_147;
  reg [31:0] dark_laplace_us_2_update_0_stage_148;
  reg [31:0] dark_laplace_us_2_update_0_stage_149;
  reg [31:0] dark_laplace_us_2_update_0_stage_150;
  reg [31:0] dark_laplace_us_2_update_0_stage_151;
  reg [31:0] dark_laplace_us_2_update_0_stage_152;
  reg [31:0] dark_laplace_us_2_update_0_stage_153;
  reg [31:0] dark_laplace_us_2_update_0_stage_154;
  reg [31:0] dark_laplace_us_2_update_0_stage_155;
  reg [31:0] dark_laplace_us_2_update_0_stage_156;
  reg [31:0] dark_laplace_us_2_update_0_stage_157;
  reg [31:0] dark_laplace_us_2_update_0_stage_158;
  reg [31:0] dark_laplace_us_2_update_0_stage_159;
  reg [31:0] dark_laplace_us_2_update_0_stage_160;
  reg [31:0] dark_laplace_us_2_update_0_stage_161;
  reg [31:0] dark_laplace_us_2_update_0_stage_162;
  reg [31:0] dark_laplace_us_2_update_0_stage_163;
  reg [31:0] dark_laplace_us_2_update_0_stage_164;
  reg [31:0] dark_laplace_us_2_update_0_stage_165;
  reg [31:0] dark_laplace_us_2_update_0_stage_166;
  reg [31:0] dark_laplace_us_2_update_0_stage_167;
  reg [31:0] dark_laplace_us_2_update_0_stage_168;
  reg [31:0] dark_laplace_us_2_update_0_stage_169;
  reg [31:0] dark_laplace_us_2_update_0_stage_170;
  reg [31:0] dark_laplace_us_2_update_0_stage_171;
  reg [31:0] dark_laplace_us_2_update_0_stage_172;
  reg [31:0] dark_laplace_us_2_update_0_stage_173;
  reg [31:0] dark_laplace_us_2_update_0_stage_174;
  reg [31:0] dark_laplace_us_2_update_0_stage_175;
  reg [31:0] dark_laplace_us_2_update_0_stage_176;
  reg [31:0] dark_laplace_us_2_update_0_stage_177;
  reg [31:0] dark_laplace_us_2_update_0_stage_178;
  reg [31:0] dark_laplace_us_2_update_0_stage_179;
  reg [31:0] dark_laplace_us_2_update_0_stage_180;
  reg [31:0] dark_laplace_us_2_update_0_stage_181;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_144;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_145;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_146;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_147;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_148;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_149;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_150;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_151;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_152;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_153;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_154;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_155;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_156;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_157;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_158;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_159;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_160;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_161;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_162;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_163;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_164;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_165;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_166;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_167;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_168;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_169;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_170;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_171;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_172;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_173;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_174;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_175;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_176;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_177;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_178;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_179;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_180;
  reg [31:0] dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_181;
  reg [31:0] final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_179;
  reg [31:0] final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_180;
  reg [31:0] final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_181;
  reg [31:0] pyramid_synthetic_exposure_fusion_update_0_stage_180;
  reg [31:0] pyramid_synthetic_exposure_fusion_update_0_stage_181;
  reg [31:0] pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127_stage_181;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_23;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_24;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_25;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_26;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_27;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_28;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_29;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_30;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_31;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_32;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_33;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_34;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_35;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_36;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_37;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_38;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_39;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_40;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_41;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_42;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_43;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_44;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_45;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_46;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_47;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_48;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_49;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_50;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_51;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_52;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_53;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_54;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_55;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_56;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_57;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_58;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_59;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_60;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_61;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_62;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_63;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_64;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_65;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_66;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_67;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_68;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_69;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_70;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_71;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_72;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_73;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_74;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_75;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_76;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_77;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_78;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_79;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_80;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_81;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_82;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_83;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_84;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_85;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_86;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_87;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_88;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_89;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_90;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_91;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_92;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_93;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_94;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_95;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_96;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_97;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_98;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_99;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_100;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_101;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_102;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_103;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_104;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_105;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_106;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_107;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_108;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_109;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_110;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_111;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_112;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_113;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_114;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_115;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_116;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_117;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_118;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_119;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_120;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_121;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_122;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_123;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_124;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_125;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_126;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_127;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_128;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_129;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_130;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_131;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_132;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_133;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_134;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_135;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_136;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_137;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_138;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_139;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_140;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_141;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_142;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_143;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_144;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_145;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_146;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_147;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_148;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_149;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_150;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_151;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_152;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_153;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_154;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_155;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_156;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_157;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_158;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_159;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_160;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_161;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_162;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_163;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_164;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_165;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_166;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_167;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_168;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_169;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_170;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_171;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_172;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_173;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_174;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_175;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_176;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_177;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_178;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_179;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_180;
  reg [31:0] dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_181;
  reg [31:0] dark_gauss_ds_1_update_0_stage_24;
  reg [31:0] dark_gauss_ds_1_update_0_stage_25;
  reg [31:0] dark_gauss_ds_1_update_0_stage_26;
  reg [31:0] dark_gauss_ds_1_update_0_stage_27;
  reg [31:0] dark_gauss_ds_1_update_0_stage_28;
  reg [31:0] dark_gauss_ds_1_update_0_stage_29;
  reg [31:0] dark_gauss_ds_1_update_0_stage_30;
  reg [31:0] dark_gauss_ds_1_update_0_stage_31;
  reg [31:0] dark_gauss_ds_1_update_0_stage_32;
  reg [31:0] dark_gauss_ds_1_update_0_stage_33;
  reg [31:0] dark_gauss_ds_1_update_0_stage_34;
  reg [31:0] dark_gauss_ds_1_update_0_stage_35;
  reg [31:0] dark_gauss_ds_1_update_0_stage_36;
  reg [31:0] dark_gauss_ds_1_update_0_stage_37;
  reg [31:0] dark_gauss_ds_1_update_0_stage_38;
  reg [31:0] dark_gauss_ds_1_update_0_stage_39;
  reg [31:0] dark_gauss_ds_1_update_0_stage_40;
  reg [31:0] dark_gauss_ds_1_update_0_stage_41;
  reg [31:0] dark_gauss_ds_1_update_0_stage_42;
  reg [31:0] dark_gauss_ds_1_update_0_stage_43;
  reg [31:0] dark_gauss_ds_1_update_0_stage_44;
  reg [31:0] dark_gauss_ds_1_update_0_stage_45;
  reg [31:0] dark_gauss_ds_1_update_0_stage_46;
  reg [31:0] dark_gauss_ds_1_update_0_stage_47;
  reg [31:0] dark_gauss_ds_1_update_0_stage_48;
  reg [31:0] dark_gauss_ds_1_update_0_stage_49;
  reg [31:0] dark_gauss_ds_1_update_0_stage_50;
  reg [31:0] dark_gauss_ds_1_update_0_stage_51;
  reg [31:0] dark_gauss_ds_1_update_0_stage_52;
  reg [31:0] dark_gauss_ds_1_update_0_stage_53;
  reg [31:0] dark_gauss_ds_1_update_0_stage_54;
  reg [31:0] dark_gauss_ds_1_update_0_stage_55;
  reg [31:0] dark_gauss_ds_1_update_0_stage_56;
  reg [31:0] dark_gauss_ds_1_update_0_stage_57;
  reg [31:0] dark_gauss_ds_1_update_0_stage_58;
  reg [31:0] dark_gauss_ds_1_update_0_stage_59;
  reg [31:0] dark_gauss_ds_1_update_0_stage_60;
  reg [31:0] dark_gauss_ds_1_update_0_stage_61;
  reg [31:0] dark_gauss_ds_1_update_0_stage_62;
  reg [31:0] dark_gauss_ds_1_update_0_stage_63;
  reg [31:0] dark_gauss_ds_1_update_0_stage_64;
  reg [31:0] dark_gauss_ds_1_update_0_stage_65;
  reg [31:0] dark_gauss_ds_1_update_0_stage_66;
  reg [31:0] dark_gauss_ds_1_update_0_stage_67;
  reg [31:0] dark_gauss_ds_1_update_0_stage_68;
  reg [31:0] dark_gauss_ds_1_update_0_stage_69;
  reg [31:0] dark_gauss_ds_1_update_0_stage_70;
  reg [31:0] dark_gauss_ds_1_update_0_stage_71;
  reg [31:0] dark_gauss_ds_1_update_0_stage_72;
  reg [31:0] dark_gauss_ds_1_update_0_stage_73;
  reg [31:0] dark_gauss_ds_1_update_0_stage_74;
  reg [31:0] dark_gauss_ds_1_update_0_stage_75;
  reg [31:0] dark_gauss_ds_1_update_0_stage_76;
  reg [31:0] dark_gauss_ds_1_update_0_stage_77;
  reg [31:0] dark_gauss_ds_1_update_0_stage_78;
  reg [31:0] dark_gauss_ds_1_update_0_stage_79;
  reg [31:0] dark_gauss_ds_1_update_0_stage_80;
  reg [31:0] dark_gauss_ds_1_update_0_stage_81;
  reg [31:0] dark_gauss_ds_1_update_0_stage_82;
  reg [31:0] dark_gauss_ds_1_update_0_stage_83;
  reg [31:0] dark_gauss_ds_1_update_0_stage_84;
  reg [31:0] dark_gauss_ds_1_update_0_stage_85;
  reg [31:0] dark_gauss_ds_1_update_0_stage_86;
  reg [31:0] dark_gauss_ds_1_update_0_stage_87;
  reg [31:0] dark_gauss_ds_1_update_0_stage_88;
  reg [31:0] dark_gauss_ds_1_update_0_stage_89;
  reg [31:0] dark_gauss_ds_1_update_0_stage_90;
  reg [31:0] dark_gauss_ds_1_update_0_stage_91;
  reg [31:0] dark_gauss_ds_1_update_0_stage_92;
  reg [31:0] dark_gauss_ds_1_update_0_stage_93;
  reg [31:0] dark_gauss_ds_1_update_0_stage_94;
  reg [31:0] dark_gauss_ds_1_update_0_stage_95;
  reg [31:0] dark_gauss_ds_1_update_0_stage_96;
  reg [31:0] dark_gauss_ds_1_update_0_stage_97;
  reg [31:0] dark_gauss_ds_1_update_0_stage_98;
  reg [31:0] dark_gauss_ds_1_update_0_stage_99;
  reg [31:0] dark_gauss_ds_1_update_0_stage_100;
  reg [31:0] dark_gauss_ds_1_update_0_stage_101;
  reg [31:0] dark_gauss_ds_1_update_0_stage_102;
  reg [31:0] dark_gauss_ds_1_update_0_stage_103;
  reg [31:0] dark_gauss_ds_1_update_0_stage_104;
  reg [31:0] dark_gauss_ds_1_update_0_stage_105;
  reg [31:0] dark_gauss_ds_1_update_0_stage_106;
  reg [31:0] dark_gauss_ds_1_update_0_stage_107;
  reg [31:0] dark_gauss_ds_1_update_0_stage_108;
  reg [31:0] dark_gauss_ds_1_update_0_stage_109;
  reg [31:0] dark_gauss_ds_1_update_0_stage_110;
  reg [31:0] dark_gauss_ds_1_update_0_stage_111;
  reg [31:0] dark_gauss_ds_1_update_0_stage_112;
  reg [31:0] dark_gauss_ds_1_update_0_stage_113;
  reg [31:0] dark_gauss_ds_1_update_0_stage_114;
  reg [31:0] dark_gauss_ds_1_update_0_stage_115;
  reg [31:0] dark_gauss_ds_1_update_0_stage_116;
  reg [31:0] dark_gauss_ds_1_update_0_stage_117;
  reg [31:0] dark_gauss_ds_1_update_0_stage_118;
  reg [31:0] dark_gauss_ds_1_update_0_stage_119;
  reg [31:0] dark_gauss_ds_1_update_0_stage_120;
  reg [31:0] dark_gauss_ds_1_update_0_stage_121;
  reg [31:0] dark_gauss_ds_1_update_0_stage_122;
  reg [31:0] dark_gauss_ds_1_update_0_stage_123;
  reg [31:0] dark_gauss_ds_1_update_0_stage_124;
  reg [31:0] dark_gauss_ds_1_update_0_stage_125;
  reg [31:0] dark_gauss_ds_1_update_0_stage_126;
  reg [31:0] dark_gauss_ds_1_update_0_stage_127;
  reg [31:0] dark_gauss_ds_1_update_0_stage_128;
  reg [31:0] dark_gauss_ds_1_update_0_stage_129;
  reg [31:0] dark_gauss_ds_1_update_0_stage_130;
  reg [31:0] dark_gauss_ds_1_update_0_stage_131;
  reg [31:0] dark_gauss_ds_1_update_0_stage_132;
  reg [31:0] dark_gauss_ds_1_update_0_stage_133;
  reg [31:0] dark_gauss_ds_1_update_0_stage_134;
  reg [31:0] dark_gauss_ds_1_update_0_stage_135;
  reg [31:0] dark_gauss_ds_1_update_0_stage_136;
  reg [31:0] dark_gauss_ds_1_update_0_stage_137;
  reg [31:0] dark_gauss_ds_1_update_0_stage_138;
  reg [31:0] dark_gauss_ds_1_update_0_stage_139;
  reg [31:0] dark_gauss_ds_1_update_0_stage_140;
  reg [31:0] dark_gauss_ds_1_update_0_stage_141;
  reg [31:0] dark_gauss_ds_1_update_0_stage_142;
  reg [31:0] dark_gauss_ds_1_update_0_stage_143;
  reg [31:0] dark_gauss_ds_1_update_0_stage_144;
  reg [31:0] dark_gauss_ds_1_update_0_stage_145;
  reg [31:0] dark_gauss_ds_1_update_0_stage_146;
  reg [31:0] dark_gauss_ds_1_update_0_stage_147;
  reg [31:0] dark_gauss_ds_1_update_0_stage_148;
  reg [31:0] dark_gauss_ds_1_update_0_stage_149;
  reg [31:0] dark_gauss_ds_1_update_0_stage_150;
  reg [31:0] dark_gauss_ds_1_update_0_stage_151;
  reg [31:0] dark_gauss_ds_1_update_0_stage_152;
  reg [31:0] dark_gauss_ds_1_update_0_stage_153;
  reg [31:0] dark_gauss_ds_1_update_0_stage_154;
  reg [31:0] dark_gauss_ds_1_update_0_stage_155;
  reg [31:0] dark_gauss_ds_1_update_0_stage_156;
  reg [31:0] dark_gauss_ds_1_update_0_stage_157;
  reg [31:0] dark_gauss_ds_1_update_0_stage_158;
  reg [31:0] dark_gauss_ds_1_update_0_stage_159;
  reg [31:0] dark_gauss_ds_1_update_0_stage_160;
  reg [31:0] dark_gauss_ds_1_update_0_stage_161;
  reg [31:0] dark_gauss_ds_1_update_0_stage_162;
  reg [31:0] dark_gauss_ds_1_update_0_stage_163;
  reg [31:0] dark_gauss_ds_1_update_0_stage_164;
  reg [31:0] dark_gauss_ds_1_update_0_stage_165;
  reg [31:0] dark_gauss_ds_1_update_0_stage_166;
  reg [31:0] dark_gauss_ds_1_update_0_stage_167;
  reg [31:0] dark_gauss_ds_1_update_0_stage_168;
  reg [31:0] dark_gauss_ds_1_update_0_stage_169;
  reg [31:0] dark_gauss_ds_1_update_0_stage_170;
  reg [31:0] dark_gauss_ds_1_update_0_stage_171;
  reg [31:0] dark_gauss_ds_1_update_0_stage_172;
  reg [31:0] dark_gauss_ds_1_update_0_stage_173;
  reg [31:0] dark_gauss_ds_1_update_0_stage_174;
  reg [31:0] dark_gauss_ds_1_update_0_stage_175;
  reg [31:0] dark_gauss_ds_1_update_0_stage_176;
  reg [31:0] dark_gauss_ds_1_update_0_stage_177;
  reg [31:0] dark_gauss_ds_1_update_0_stage_178;
  reg [31:0] dark_gauss_ds_1_update_0_stage_179;
  reg [31:0] dark_gauss_ds_1_update_0_stage_180;
  reg [31:0] dark_gauss_ds_1_update_0_stage_181;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_25;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_26;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_27;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_28;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_29;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_30;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_31;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_32;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_33;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_34;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_35;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_36;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_37;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_38;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_39;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_40;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_41;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_42;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_43;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_44;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_45;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_46;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_47;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_48;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_49;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_50;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_51;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_52;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_53;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_54;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_55;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_56;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_57;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_58;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_59;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_60;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_61;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_62;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_63;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_64;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_65;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_66;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_67;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_68;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_69;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_70;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_71;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_72;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_73;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_74;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_75;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_76;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_77;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_78;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_79;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_80;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_81;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_82;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_83;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_84;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_85;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_86;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_87;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_88;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_89;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_90;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_91;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_92;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_93;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_94;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_95;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_96;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_97;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_98;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_99;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_100;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_101;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_102;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_103;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_104;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_105;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_106;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_107;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_108;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_109;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_110;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_111;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_112;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_113;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_114;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_115;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_116;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_117;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_118;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_119;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_120;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_121;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_122;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_123;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_124;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_125;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_126;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_127;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_128;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_129;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_130;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_131;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_132;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_133;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_134;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_135;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_136;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_137;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_138;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_139;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_140;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_141;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_142;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_143;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_144;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_145;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_146;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_147;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_148;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_149;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_150;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_151;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_152;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_153;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_154;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_155;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_156;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_157;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_158;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_159;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_160;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_161;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_162;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_163;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_164;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_165;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_166;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_167;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_168;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_169;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_170;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_171;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_172;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_173;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_174;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_175;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_176;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_177;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_178;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_179;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_180;
  reg [31:0] dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_181;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_31;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_32;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_33;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_34;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_35;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_36;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_37;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_38;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_39;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_40;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_41;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_42;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_43;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_44;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_45;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_46;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_47;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_48;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_49;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_50;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_51;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_52;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_53;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_54;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_55;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_56;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_57;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_58;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_59;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_60;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_61;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_62;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_63;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_64;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_65;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_66;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_67;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_68;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_69;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_70;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_71;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_72;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_73;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_74;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_75;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_76;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_77;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_78;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_79;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_80;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_81;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_82;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_83;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_84;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_85;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_86;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_87;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_88;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_89;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_90;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_91;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_92;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_93;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_94;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_95;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_96;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_97;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_98;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_99;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_100;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_101;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_102;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_103;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_104;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_105;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_106;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_107;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_108;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_109;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_110;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_111;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_112;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_113;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_114;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_115;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_116;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_117;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_118;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_119;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_120;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_121;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_122;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_123;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_124;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_125;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_126;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_127;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_128;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_129;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_130;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_131;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_132;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_133;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_134;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_135;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_136;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_137;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_138;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_139;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_140;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_141;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_142;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_143;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_144;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_145;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_146;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_147;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_148;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_149;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_150;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_151;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_152;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_153;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_154;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_155;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_156;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_157;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_158;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_159;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_160;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_161;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_162;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_163;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_164;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_165;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_166;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_167;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_168;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_169;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_170;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_171;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_172;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_173;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_174;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_175;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_176;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_177;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_178;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_179;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_180;
  reg [31:0] dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_181;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_32;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_33;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_34;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_35;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_36;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_37;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_38;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_39;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_40;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_41;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_42;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_43;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_44;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_45;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_46;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_47;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_48;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_49;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_50;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_51;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_52;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_53;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_54;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_55;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_56;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_57;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_58;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_59;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_60;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_61;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_62;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_63;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_64;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_65;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_66;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_67;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_68;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_69;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_70;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_71;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_72;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_73;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_74;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_75;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_76;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_77;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_78;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_79;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_80;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_81;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_82;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_83;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_84;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_85;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_86;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_87;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_88;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_89;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_90;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_91;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_92;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_93;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_94;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_95;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_96;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_97;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_98;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_99;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_100;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_101;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_102;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_103;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_104;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_105;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_106;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_107;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_108;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_109;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_110;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_111;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_112;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_113;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_114;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_115;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_116;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_117;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_118;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_119;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_120;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_121;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_122;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_123;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_124;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_125;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_126;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_127;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_128;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_129;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_130;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_131;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_132;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_133;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_134;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_135;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_136;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_137;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_138;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_139;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_140;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_141;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_142;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_143;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_144;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_145;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_146;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_147;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_148;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_149;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_150;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_151;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_152;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_153;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_154;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_155;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_156;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_157;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_158;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_159;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_160;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_161;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_162;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_163;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_164;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_165;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_166;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_167;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_168;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_169;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_170;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_171;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_172;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_173;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_174;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_175;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_176;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_177;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_178;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_179;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_180;
  reg [31:0] bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_181;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_29;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_30;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_31;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_32;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_33;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_34;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_35;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_36;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_37;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_38;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_39;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_40;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_41;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_42;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_43;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_44;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_45;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_46;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_47;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_48;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_49;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_50;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_51;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_52;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_53;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_54;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_55;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_56;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_57;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_58;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_59;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_60;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_61;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_62;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_63;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_64;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_65;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_66;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_67;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_68;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_69;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_70;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_71;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_72;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_73;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_74;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_75;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_76;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_77;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_78;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_79;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_80;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_81;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_82;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_83;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_84;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_85;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_86;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_87;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_88;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_89;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_90;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_91;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_92;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_93;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_94;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_95;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_96;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_97;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_98;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_99;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_100;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_101;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_102;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_103;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_104;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_105;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_106;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_107;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_108;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_109;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_110;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_111;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_112;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_113;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_114;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_115;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_116;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_117;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_118;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_119;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_120;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_121;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_122;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_123;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_124;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_125;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_126;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_127;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_128;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_129;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_130;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_131;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_132;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_133;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_134;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_135;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_136;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_137;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_138;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_139;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_140;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_141;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_142;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_143;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_144;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_145;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_146;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_147;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_148;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_149;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_150;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_151;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_152;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_153;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_154;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_155;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_156;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_157;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_158;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_159;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_160;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_161;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_162;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_163;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_164;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_165;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_166;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_167;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_168;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_169;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_170;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_171;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_172;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_173;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_174;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_175;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_176;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_177;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_178;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_179;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_180;
  reg [287:0] dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_181;
  reg [31:0] dark_gauss_blur_2_update_0_stage_30;
  reg [31:0] dark_gauss_blur_2_update_0_stage_31;
  reg [31:0] dark_gauss_blur_2_update_0_stage_32;
  reg [31:0] dark_gauss_blur_2_update_0_stage_33;
  reg [31:0] dark_gauss_blur_2_update_0_stage_34;
  reg [31:0] dark_gauss_blur_2_update_0_stage_35;
  reg [31:0] dark_gauss_blur_2_update_0_stage_36;
  reg [31:0] dark_gauss_blur_2_update_0_stage_37;
  reg [31:0] dark_gauss_blur_2_update_0_stage_38;
  reg [31:0] dark_gauss_blur_2_update_0_stage_39;
  reg [31:0] dark_gauss_blur_2_update_0_stage_40;
  reg [31:0] dark_gauss_blur_2_update_0_stage_41;
  reg [31:0] dark_gauss_blur_2_update_0_stage_42;
  reg [31:0] dark_gauss_blur_2_update_0_stage_43;
  reg [31:0] dark_gauss_blur_2_update_0_stage_44;
  reg [31:0] dark_gauss_blur_2_update_0_stage_45;
  reg [31:0] dark_gauss_blur_2_update_0_stage_46;
  reg [31:0] dark_gauss_blur_2_update_0_stage_47;
  reg [31:0] dark_gauss_blur_2_update_0_stage_48;
  reg [31:0] dark_gauss_blur_2_update_0_stage_49;
  reg [31:0] dark_gauss_blur_2_update_0_stage_50;
  reg [31:0] dark_gauss_blur_2_update_0_stage_51;
  reg [31:0] dark_gauss_blur_2_update_0_stage_52;
  reg [31:0] dark_gauss_blur_2_update_0_stage_53;
  reg [31:0] dark_gauss_blur_2_update_0_stage_54;
  reg [31:0] dark_gauss_blur_2_update_0_stage_55;
  reg [31:0] dark_gauss_blur_2_update_0_stage_56;
  reg [31:0] dark_gauss_blur_2_update_0_stage_57;
  reg [31:0] dark_gauss_blur_2_update_0_stage_58;
  reg [31:0] dark_gauss_blur_2_update_0_stage_59;
  reg [31:0] dark_gauss_blur_2_update_0_stage_60;
  reg [31:0] dark_gauss_blur_2_update_0_stage_61;
  reg [31:0] dark_gauss_blur_2_update_0_stage_62;
  reg [31:0] dark_gauss_blur_2_update_0_stage_63;
  reg [31:0] dark_gauss_blur_2_update_0_stage_64;
  reg [31:0] dark_gauss_blur_2_update_0_stage_65;
  reg [31:0] dark_gauss_blur_2_update_0_stage_66;
  reg [31:0] dark_gauss_blur_2_update_0_stage_67;
  reg [31:0] dark_gauss_blur_2_update_0_stage_68;
  reg [31:0] dark_gauss_blur_2_update_0_stage_69;
  reg [31:0] dark_gauss_blur_2_update_0_stage_70;
  reg [31:0] dark_gauss_blur_2_update_0_stage_71;
  reg [31:0] dark_gauss_blur_2_update_0_stage_72;
  reg [31:0] dark_gauss_blur_2_update_0_stage_73;
  reg [31:0] dark_gauss_blur_2_update_0_stage_74;
  reg [31:0] dark_gauss_blur_2_update_0_stage_75;
  reg [31:0] dark_gauss_blur_2_update_0_stage_76;
  reg [31:0] dark_gauss_blur_2_update_0_stage_77;
  reg [31:0] dark_gauss_blur_2_update_0_stage_78;
  reg [31:0] dark_gauss_blur_2_update_0_stage_79;
  reg [31:0] dark_gauss_blur_2_update_0_stage_80;
  reg [31:0] dark_gauss_blur_2_update_0_stage_81;
  reg [31:0] dark_gauss_blur_2_update_0_stage_82;
  reg [31:0] dark_gauss_blur_2_update_0_stage_83;
  reg [31:0] dark_gauss_blur_2_update_0_stage_84;
  reg [31:0] dark_gauss_blur_2_update_0_stage_85;
  reg [31:0] dark_gauss_blur_2_update_0_stage_86;
  reg [31:0] dark_gauss_blur_2_update_0_stage_87;
  reg [31:0] dark_gauss_blur_2_update_0_stage_88;
  reg [31:0] dark_gauss_blur_2_update_0_stage_89;
  reg [31:0] dark_gauss_blur_2_update_0_stage_90;
  reg [31:0] dark_gauss_blur_2_update_0_stage_91;
  reg [31:0] dark_gauss_blur_2_update_0_stage_92;
  reg [31:0] dark_gauss_blur_2_update_0_stage_93;
  reg [31:0] dark_gauss_blur_2_update_0_stage_94;
  reg [31:0] dark_gauss_blur_2_update_0_stage_95;
  reg [31:0] dark_gauss_blur_2_update_0_stage_96;
  reg [31:0] dark_gauss_blur_2_update_0_stage_97;
  reg [31:0] dark_gauss_blur_2_update_0_stage_98;
  reg [31:0] dark_gauss_blur_2_update_0_stage_99;
  reg [31:0] dark_gauss_blur_2_update_0_stage_100;
  reg [31:0] dark_gauss_blur_2_update_0_stage_101;
  reg [31:0] dark_gauss_blur_2_update_0_stage_102;
  reg [31:0] dark_gauss_blur_2_update_0_stage_103;
  reg [31:0] dark_gauss_blur_2_update_0_stage_104;
  reg [31:0] dark_gauss_blur_2_update_0_stage_105;
  reg [31:0] dark_gauss_blur_2_update_0_stage_106;
  reg [31:0] dark_gauss_blur_2_update_0_stage_107;
  reg [31:0] dark_gauss_blur_2_update_0_stage_108;
  reg [31:0] dark_gauss_blur_2_update_0_stage_109;
  reg [31:0] dark_gauss_blur_2_update_0_stage_110;
  reg [31:0] dark_gauss_blur_2_update_0_stage_111;
  reg [31:0] dark_gauss_blur_2_update_0_stage_112;
  reg [31:0] dark_gauss_blur_2_update_0_stage_113;
  reg [31:0] dark_gauss_blur_2_update_0_stage_114;
  reg [31:0] dark_gauss_blur_2_update_0_stage_115;
  reg [31:0] dark_gauss_blur_2_update_0_stage_116;
  reg [31:0] dark_gauss_blur_2_update_0_stage_117;
  reg [31:0] dark_gauss_blur_2_update_0_stage_118;
  reg [31:0] dark_gauss_blur_2_update_0_stage_119;
  reg [31:0] dark_gauss_blur_2_update_0_stage_120;
  reg [31:0] dark_gauss_blur_2_update_0_stage_121;
  reg [31:0] dark_gauss_blur_2_update_0_stage_122;
  reg [31:0] dark_gauss_blur_2_update_0_stage_123;
  reg [31:0] dark_gauss_blur_2_update_0_stage_124;
  reg [31:0] dark_gauss_blur_2_update_0_stage_125;
  reg [31:0] dark_gauss_blur_2_update_0_stage_126;
  reg [31:0] dark_gauss_blur_2_update_0_stage_127;
  reg [31:0] dark_gauss_blur_2_update_0_stage_128;
  reg [31:0] dark_gauss_blur_2_update_0_stage_129;
  reg [31:0] dark_gauss_blur_2_update_0_stage_130;
  reg [31:0] dark_gauss_blur_2_update_0_stage_131;
  reg [31:0] dark_gauss_blur_2_update_0_stage_132;
  reg [31:0] dark_gauss_blur_2_update_0_stage_133;
  reg [31:0] dark_gauss_blur_2_update_0_stage_134;
  reg [31:0] dark_gauss_blur_2_update_0_stage_135;
  reg [31:0] dark_gauss_blur_2_update_0_stage_136;
  reg [31:0] dark_gauss_blur_2_update_0_stage_137;
  reg [31:0] dark_gauss_blur_2_update_0_stage_138;
  reg [31:0] dark_gauss_blur_2_update_0_stage_139;
  reg [31:0] dark_gauss_blur_2_update_0_stage_140;
  reg [31:0] dark_gauss_blur_2_update_0_stage_141;
  reg [31:0] dark_gauss_blur_2_update_0_stage_142;
  reg [31:0] dark_gauss_blur_2_update_0_stage_143;
  reg [31:0] dark_gauss_blur_2_update_0_stage_144;
  reg [31:0] dark_gauss_blur_2_update_0_stage_145;
  reg [31:0] dark_gauss_blur_2_update_0_stage_146;
  reg [31:0] dark_gauss_blur_2_update_0_stage_147;
  reg [31:0] dark_gauss_blur_2_update_0_stage_148;
  reg [31:0] dark_gauss_blur_2_update_0_stage_149;
  reg [31:0] dark_gauss_blur_2_update_0_stage_150;
  reg [31:0] dark_gauss_blur_2_update_0_stage_151;
  reg [31:0] dark_gauss_blur_2_update_0_stage_152;
  reg [31:0] dark_gauss_blur_2_update_0_stage_153;
  reg [31:0] dark_gauss_blur_2_update_0_stage_154;
  reg [31:0] dark_gauss_blur_2_update_0_stage_155;
  reg [31:0] dark_gauss_blur_2_update_0_stage_156;
  reg [31:0] dark_gauss_blur_2_update_0_stage_157;
  reg [31:0] dark_gauss_blur_2_update_0_stage_158;
  reg [31:0] dark_gauss_blur_2_update_0_stage_159;
  reg [31:0] dark_gauss_blur_2_update_0_stage_160;
  reg [31:0] dark_gauss_blur_2_update_0_stage_161;
  reg [31:0] dark_gauss_blur_2_update_0_stage_162;
  reg [31:0] dark_gauss_blur_2_update_0_stage_163;
  reg [31:0] dark_gauss_blur_2_update_0_stage_164;
  reg [31:0] dark_gauss_blur_2_update_0_stage_165;
  reg [31:0] dark_gauss_blur_2_update_0_stage_166;
  reg [31:0] dark_gauss_blur_2_update_0_stage_167;
  reg [31:0] dark_gauss_blur_2_update_0_stage_168;
  reg [31:0] dark_gauss_blur_2_update_0_stage_169;
  reg [31:0] dark_gauss_blur_2_update_0_stage_170;
  reg [31:0] dark_gauss_blur_2_update_0_stage_171;
  reg [31:0] dark_gauss_blur_2_update_0_stage_172;
  reg [31:0] dark_gauss_blur_2_update_0_stage_173;
  reg [31:0] dark_gauss_blur_2_update_0_stage_174;
  reg [31:0] dark_gauss_blur_2_update_0_stage_175;
  reg [31:0] dark_gauss_blur_2_update_0_stage_176;
  reg [31:0] dark_gauss_blur_2_update_0_stage_177;
  reg [31:0] dark_gauss_blur_2_update_0_stage_178;
  reg [31:0] dark_gauss_blur_2_update_0_stage_179;
  reg [31:0] dark_gauss_blur_2_update_0_stage_180;
  reg [31:0] dark_gauss_blur_2_update_0_stage_181;
  reg [31:0] bright_gauss_ds_1_update_0_stage_33;
  reg [31:0] bright_gauss_ds_1_update_0_stage_34;
  reg [31:0] bright_gauss_ds_1_update_0_stage_35;
  reg [31:0] bright_gauss_ds_1_update_0_stage_36;
  reg [31:0] bright_gauss_ds_1_update_0_stage_37;
  reg [31:0] bright_gauss_ds_1_update_0_stage_38;
  reg [31:0] bright_gauss_ds_1_update_0_stage_39;
  reg [31:0] bright_gauss_ds_1_update_0_stage_40;
  reg [31:0] bright_gauss_ds_1_update_0_stage_41;
  reg [31:0] bright_gauss_ds_1_update_0_stage_42;
  reg [31:0] bright_gauss_ds_1_update_0_stage_43;
  reg [31:0] bright_gauss_ds_1_update_0_stage_44;
  reg [31:0] bright_gauss_ds_1_update_0_stage_45;
  reg [31:0] bright_gauss_ds_1_update_0_stage_46;
  reg [31:0] bright_gauss_ds_1_update_0_stage_47;
  reg [31:0] bright_gauss_ds_1_update_0_stage_48;
  reg [31:0] bright_gauss_ds_1_update_0_stage_49;
  reg [31:0] bright_gauss_ds_1_update_0_stage_50;
  reg [31:0] bright_gauss_ds_1_update_0_stage_51;
  reg [31:0] bright_gauss_ds_1_update_0_stage_52;
  reg [31:0] bright_gauss_ds_1_update_0_stage_53;
  reg [31:0] bright_gauss_ds_1_update_0_stage_54;
  reg [31:0] bright_gauss_ds_1_update_0_stage_55;
  reg [31:0] bright_gauss_ds_1_update_0_stage_56;
  reg [31:0] bright_gauss_ds_1_update_0_stage_57;
  reg [31:0] bright_gauss_ds_1_update_0_stage_58;
  reg [31:0] bright_gauss_ds_1_update_0_stage_59;
  reg [31:0] bright_gauss_ds_1_update_0_stage_60;
  reg [31:0] bright_gauss_ds_1_update_0_stage_61;
  reg [31:0] bright_gauss_ds_1_update_0_stage_62;
  reg [31:0] bright_gauss_ds_1_update_0_stage_63;
  reg [31:0] bright_gauss_ds_1_update_0_stage_64;
  reg [31:0] bright_gauss_ds_1_update_0_stage_65;
  reg [31:0] bright_gauss_ds_1_update_0_stage_66;
  reg [31:0] bright_gauss_ds_1_update_0_stage_67;
  reg [31:0] bright_gauss_ds_1_update_0_stage_68;
  reg [31:0] bright_gauss_ds_1_update_0_stage_69;
  reg [31:0] bright_gauss_ds_1_update_0_stage_70;
  reg [31:0] bright_gauss_ds_1_update_0_stage_71;
  reg [31:0] bright_gauss_ds_1_update_0_stage_72;
  reg [31:0] bright_gauss_ds_1_update_0_stage_73;
  reg [31:0] bright_gauss_ds_1_update_0_stage_74;
  reg [31:0] bright_gauss_ds_1_update_0_stage_75;
  reg [31:0] bright_gauss_ds_1_update_0_stage_76;
  reg [31:0] bright_gauss_ds_1_update_0_stage_77;
  reg [31:0] bright_gauss_ds_1_update_0_stage_78;
  reg [31:0] bright_gauss_ds_1_update_0_stage_79;
  reg [31:0] bright_gauss_ds_1_update_0_stage_80;
  reg [31:0] bright_gauss_ds_1_update_0_stage_81;
  reg [31:0] bright_gauss_ds_1_update_0_stage_82;
  reg [31:0] bright_gauss_ds_1_update_0_stage_83;
  reg [31:0] bright_gauss_ds_1_update_0_stage_84;
  reg [31:0] bright_gauss_ds_1_update_0_stage_85;
  reg [31:0] bright_gauss_ds_1_update_0_stage_86;
  reg [31:0] bright_gauss_ds_1_update_0_stage_87;
  reg [31:0] bright_gauss_ds_1_update_0_stage_88;
  reg [31:0] bright_gauss_ds_1_update_0_stage_89;
  reg [31:0] bright_gauss_ds_1_update_0_stage_90;
  reg [31:0] bright_gauss_ds_1_update_0_stage_91;
  reg [31:0] bright_gauss_ds_1_update_0_stage_92;
  reg [31:0] bright_gauss_ds_1_update_0_stage_93;
  reg [31:0] bright_gauss_ds_1_update_0_stage_94;
  reg [31:0] bright_gauss_ds_1_update_0_stage_95;
  reg [31:0] bright_gauss_ds_1_update_0_stage_96;
  reg [31:0] bright_gauss_ds_1_update_0_stage_97;
  reg [31:0] bright_gauss_ds_1_update_0_stage_98;
  reg [31:0] bright_gauss_ds_1_update_0_stage_99;
  reg [31:0] bright_gauss_ds_1_update_0_stage_100;
  reg [31:0] bright_gauss_ds_1_update_0_stage_101;
  reg [31:0] bright_gauss_ds_1_update_0_stage_102;
  reg [31:0] bright_gauss_ds_1_update_0_stage_103;
  reg [31:0] bright_gauss_ds_1_update_0_stage_104;
  reg [31:0] bright_gauss_ds_1_update_0_stage_105;
  reg [31:0] bright_gauss_ds_1_update_0_stage_106;
  reg [31:0] bright_gauss_ds_1_update_0_stage_107;
  reg [31:0] bright_gauss_ds_1_update_0_stage_108;
  reg [31:0] bright_gauss_ds_1_update_0_stage_109;
  reg [31:0] bright_gauss_ds_1_update_0_stage_110;
  reg [31:0] bright_gauss_ds_1_update_0_stage_111;
  reg [31:0] bright_gauss_ds_1_update_0_stage_112;
  reg [31:0] bright_gauss_ds_1_update_0_stage_113;
  reg [31:0] bright_gauss_ds_1_update_0_stage_114;
  reg [31:0] bright_gauss_ds_1_update_0_stage_115;
  reg [31:0] bright_gauss_ds_1_update_0_stage_116;
  reg [31:0] bright_gauss_ds_1_update_0_stage_117;
  reg [31:0] bright_gauss_ds_1_update_0_stage_118;
  reg [31:0] bright_gauss_ds_1_update_0_stage_119;
  reg [31:0] bright_gauss_ds_1_update_0_stage_120;
  reg [31:0] bright_gauss_ds_1_update_0_stage_121;
  reg [31:0] bright_gauss_ds_1_update_0_stage_122;
  reg [31:0] bright_gauss_ds_1_update_0_stage_123;
  reg [31:0] bright_gauss_ds_1_update_0_stage_124;
  reg [31:0] bright_gauss_ds_1_update_0_stage_125;
  reg [31:0] bright_gauss_ds_1_update_0_stage_126;
  reg [31:0] bright_gauss_ds_1_update_0_stage_127;
  reg [31:0] bright_gauss_ds_1_update_0_stage_128;
  reg [31:0] bright_gauss_ds_1_update_0_stage_129;
  reg [31:0] bright_gauss_ds_1_update_0_stage_130;
  reg [31:0] bright_gauss_ds_1_update_0_stage_131;
  reg [31:0] bright_gauss_ds_1_update_0_stage_132;
  reg [31:0] bright_gauss_ds_1_update_0_stage_133;
  reg [31:0] bright_gauss_ds_1_update_0_stage_134;
  reg [31:0] bright_gauss_ds_1_update_0_stage_135;
  reg [31:0] bright_gauss_ds_1_update_0_stage_136;
  reg [31:0] bright_gauss_ds_1_update_0_stage_137;
  reg [31:0] bright_gauss_ds_1_update_0_stage_138;
  reg [31:0] bright_gauss_ds_1_update_0_stage_139;
  reg [31:0] bright_gauss_ds_1_update_0_stage_140;
  reg [31:0] bright_gauss_ds_1_update_0_stage_141;
  reg [31:0] bright_gauss_ds_1_update_0_stage_142;
  reg [31:0] bright_gauss_ds_1_update_0_stage_143;
  reg [31:0] bright_gauss_ds_1_update_0_stage_144;
  reg [31:0] bright_gauss_ds_1_update_0_stage_145;
  reg [31:0] bright_gauss_ds_1_update_0_stage_146;
  reg [31:0] bright_gauss_ds_1_update_0_stage_147;
  reg [31:0] bright_gauss_ds_1_update_0_stage_148;
  reg [31:0] bright_gauss_ds_1_update_0_stage_149;
  reg [31:0] bright_gauss_ds_1_update_0_stage_150;
  reg [31:0] bright_gauss_ds_1_update_0_stage_151;
  reg [31:0] bright_gauss_ds_1_update_0_stage_152;
  reg [31:0] bright_gauss_ds_1_update_0_stage_153;
  reg [31:0] bright_gauss_ds_1_update_0_stage_154;
  reg [31:0] bright_gauss_ds_1_update_0_stage_155;
  reg [31:0] bright_gauss_ds_1_update_0_stage_156;
  reg [31:0] bright_gauss_ds_1_update_0_stage_157;
  reg [31:0] bright_gauss_ds_1_update_0_stage_158;
  reg [31:0] bright_gauss_ds_1_update_0_stage_159;
  reg [31:0] bright_gauss_ds_1_update_0_stage_160;
  reg [31:0] bright_gauss_ds_1_update_0_stage_161;
  reg [31:0] bright_gauss_ds_1_update_0_stage_162;
  reg [31:0] bright_gauss_ds_1_update_0_stage_163;
  reg [31:0] bright_gauss_ds_1_update_0_stage_164;
  reg [31:0] bright_gauss_ds_1_update_0_stage_165;
  reg [31:0] bright_gauss_ds_1_update_0_stage_166;
  reg [31:0] bright_gauss_ds_1_update_0_stage_167;
  reg [31:0] bright_gauss_ds_1_update_0_stage_168;
  reg [31:0] bright_gauss_ds_1_update_0_stage_169;
  reg [31:0] bright_gauss_ds_1_update_0_stage_170;
  reg [31:0] bright_gauss_ds_1_update_0_stage_171;
  reg [31:0] bright_gauss_ds_1_update_0_stage_172;
  reg [31:0] bright_gauss_ds_1_update_0_stage_173;
  reg [31:0] bright_gauss_ds_1_update_0_stage_174;
  reg [31:0] bright_gauss_ds_1_update_0_stage_175;
  reg [31:0] bright_gauss_ds_1_update_0_stage_176;
  reg [31:0] bright_gauss_ds_1_update_0_stage_177;
  reg [31:0] bright_gauss_ds_1_update_0_stage_178;
  reg [31:0] bright_gauss_ds_1_update_0_stage_179;
  reg [31:0] bright_gauss_ds_1_update_0_stage_180;
  reg [31:0] bright_gauss_ds_1_update_0_stage_181;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_34;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_35;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_36;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_37;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_38;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_39;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_40;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_41;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_42;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_43;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_44;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_45;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_46;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_47;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_48;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_49;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_50;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_51;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_52;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_53;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_54;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_55;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_56;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_57;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_58;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_59;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_60;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_61;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_62;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_63;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_64;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_65;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_66;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_67;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_68;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_69;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_70;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_71;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_72;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_73;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_74;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_75;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_76;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_77;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_78;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_79;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_80;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_81;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_82;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_83;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_84;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_85;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_86;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_87;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_88;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_89;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_90;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_91;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_92;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_93;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_94;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_95;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_96;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_97;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_98;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_99;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_100;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_101;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_102;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_103;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_104;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_105;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_106;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_107;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_108;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_109;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_110;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_111;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_112;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_113;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_114;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_115;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_116;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_117;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_118;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_119;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_120;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_121;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_122;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_123;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_124;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_125;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_126;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_127;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_128;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_129;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_130;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_131;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_132;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_133;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_134;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_135;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_136;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_137;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_138;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_139;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_140;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_141;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_142;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_143;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_144;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_145;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_146;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_147;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_148;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_149;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_150;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_151;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_152;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_153;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_154;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_155;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_156;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_157;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_158;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_159;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_160;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_161;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_162;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_163;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_164;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_165;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_166;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_167;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_168;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_169;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_170;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_171;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_172;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_173;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_174;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_175;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_176;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_177;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_178;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_179;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_180;
  reg [31:0] bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_181;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_69;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_70;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_71;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_72;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_73;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_74;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_75;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_76;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_77;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_78;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_79;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_80;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_81;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_82;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_83;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_84;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_85;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_86;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_87;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_88;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_89;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_90;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_91;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_92;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_93;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_94;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_95;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_96;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_97;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_98;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_99;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_100;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_101;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_102;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_103;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_104;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_105;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_106;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_107;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_108;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_109;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_110;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_111;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_112;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_113;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_114;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_115;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_116;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_117;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_118;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_119;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_120;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_121;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_122;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_123;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_124;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_125;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_126;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_127;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_128;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_129;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_130;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_131;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_132;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_133;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_134;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_135;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_136;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_137;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_138;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_139;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_140;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_141;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_142;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_143;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_144;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_145;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_146;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_147;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_148;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_149;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_150;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_151;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_152;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_153;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_154;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_155;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_156;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_157;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_158;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_159;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_160;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_161;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_162;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_163;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_164;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_165;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_166;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_167;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_168;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_169;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_170;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_171;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_172;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_173;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_174;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_175;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_176;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_177;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_178;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_179;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_180;
  reg [31:0] weight_sums_dark_weights_normed_update_0_read_read_46_stage_181;
  reg [31:0] dark_weights_normed_update_0_stage_70;
  reg [31:0] dark_weights_normed_update_0_stage_71;
  reg [31:0] dark_weights_normed_update_0_stage_72;
  reg [31:0] dark_weights_normed_update_0_stage_73;
  reg [31:0] dark_weights_normed_update_0_stage_74;
  reg [31:0] dark_weights_normed_update_0_stage_75;
  reg [31:0] dark_weights_normed_update_0_stage_76;
  reg [31:0] dark_weights_normed_update_0_stage_77;
  reg [31:0] dark_weights_normed_update_0_stage_78;
  reg [31:0] dark_weights_normed_update_0_stage_79;
  reg [31:0] dark_weights_normed_update_0_stage_80;
  reg [31:0] dark_weights_normed_update_0_stage_81;
  reg [31:0] dark_weights_normed_update_0_stage_82;
  reg [31:0] dark_weights_normed_update_0_stage_83;
  reg [31:0] dark_weights_normed_update_0_stage_84;
  reg [31:0] dark_weights_normed_update_0_stage_85;
  reg [31:0] dark_weights_normed_update_0_stage_86;
  reg [31:0] dark_weights_normed_update_0_stage_87;
  reg [31:0] dark_weights_normed_update_0_stage_88;
  reg [31:0] dark_weights_normed_update_0_stage_89;
  reg [31:0] dark_weights_normed_update_0_stage_90;
  reg [31:0] dark_weights_normed_update_0_stage_91;
  reg [31:0] dark_weights_normed_update_0_stage_92;
  reg [31:0] dark_weights_normed_update_0_stage_93;
  reg [31:0] dark_weights_normed_update_0_stage_94;
  reg [31:0] dark_weights_normed_update_0_stage_95;
  reg [31:0] dark_weights_normed_update_0_stage_96;
  reg [31:0] dark_weights_normed_update_0_stage_97;
  reg [31:0] dark_weights_normed_update_0_stage_98;
  reg [31:0] dark_weights_normed_update_0_stage_99;
  reg [31:0] dark_weights_normed_update_0_stage_100;
  reg [31:0] dark_weights_normed_update_0_stage_101;
  reg [31:0] dark_weights_normed_update_0_stage_102;
  reg [31:0] dark_weights_normed_update_0_stage_103;
  reg [31:0] dark_weights_normed_update_0_stage_104;
  reg [31:0] dark_weights_normed_update_0_stage_105;
  reg [31:0] dark_weights_normed_update_0_stage_106;
  reg [31:0] dark_weights_normed_update_0_stage_107;
  reg [31:0] dark_weights_normed_update_0_stage_108;
  reg [31:0] dark_weights_normed_update_0_stage_109;
  reg [31:0] dark_weights_normed_update_0_stage_110;
  reg [31:0] dark_weights_normed_update_0_stage_111;
  reg [31:0] dark_weights_normed_update_0_stage_112;
  reg [31:0] dark_weights_normed_update_0_stage_113;
  reg [31:0] dark_weights_normed_update_0_stage_114;
  reg [31:0] dark_weights_normed_update_0_stage_115;
  reg [31:0] dark_weights_normed_update_0_stage_116;
  reg [31:0] dark_weights_normed_update_0_stage_117;
  reg [31:0] dark_weights_normed_update_0_stage_118;
  reg [31:0] dark_weights_normed_update_0_stage_119;
  reg [31:0] dark_weights_normed_update_0_stage_120;
  reg [31:0] dark_weights_normed_update_0_stage_121;
  reg [31:0] dark_weights_normed_update_0_stage_122;
  reg [31:0] dark_weights_normed_update_0_stage_123;
  reg [31:0] dark_weights_normed_update_0_stage_124;
  reg [31:0] dark_weights_normed_update_0_stage_125;
  reg [31:0] dark_weights_normed_update_0_stage_126;
  reg [31:0] dark_weights_normed_update_0_stage_127;
  reg [31:0] dark_weights_normed_update_0_stage_128;
  reg [31:0] dark_weights_normed_update_0_stage_129;
  reg [31:0] dark_weights_normed_update_0_stage_130;
  reg [31:0] dark_weights_normed_update_0_stage_131;
  reg [31:0] dark_weights_normed_update_0_stage_132;
  reg [31:0] dark_weights_normed_update_0_stage_133;
  reg [31:0] dark_weights_normed_update_0_stage_134;
  reg [31:0] dark_weights_normed_update_0_stage_135;
  reg [31:0] dark_weights_normed_update_0_stage_136;
  reg [31:0] dark_weights_normed_update_0_stage_137;
  reg [31:0] dark_weights_normed_update_0_stage_138;
  reg [31:0] dark_weights_normed_update_0_stage_139;
  reg [31:0] dark_weights_normed_update_0_stage_140;
  reg [31:0] dark_weights_normed_update_0_stage_141;
  reg [31:0] dark_weights_normed_update_0_stage_142;
  reg [31:0] dark_weights_normed_update_0_stage_143;
  reg [31:0] dark_weights_normed_update_0_stage_144;
  reg [31:0] dark_weights_normed_update_0_stage_145;
  reg [31:0] dark_weights_normed_update_0_stage_146;
  reg [31:0] dark_weights_normed_update_0_stage_147;
  reg [31:0] dark_weights_normed_update_0_stage_148;
  reg [31:0] dark_weights_normed_update_0_stage_149;
  reg [31:0] dark_weights_normed_update_0_stage_150;
  reg [31:0] dark_weights_normed_update_0_stage_151;
  reg [31:0] dark_weights_normed_update_0_stage_152;
  reg [31:0] dark_weights_normed_update_0_stage_153;
  reg [31:0] dark_weights_normed_update_0_stage_154;
  reg [31:0] dark_weights_normed_update_0_stage_155;
  reg [31:0] dark_weights_normed_update_0_stage_156;
  reg [31:0] dark_weights_normed_update_0_stage_157;
  reg [31:0] dark_weights_normed_update_0_stage_158;
  reg [31:0] dark_weights_normed_update_0_stage_159;
  reg [31:0] dark_weights_normed_update_0_stage_160;
  reg [31:0] dark_weights_normed_update_0_stage_161;
  reg [31:0] dark_weights_normed_update_0_stage_162;
  reg [31:0] dark_weights_normed_update_0_stage_163;
  reg [31:0] dark_weights_normed_update_0_stage_164;
  reg [31:0] dark_weights_normed_update_0_stage_165;
  reg [31:0] dark_weights_normed_update_0_stage_166;
  reg [31:0] dark_weights_normed_update_0_stage_167;
  reg [31:0] dark_weights_normed_update_0_stage_168;
  reg [31:0] dark_weights_normed_update_0_stage_169;
  reg [31:0] dark_weights_normed_update_0_stage_170;
  reg [31:0] dark_weights_normed_update_0_stage_171;
  reg [31:0] dark_weights_normed_update_0_stage_172;
  reg [31:0] dark_weights_normed_update_0_stage_173;
  reg [31:0] dark_weights_normed_update_0_stage_174;
  reg [31:0] dark_weights_normed_update_0_stage_175;
  reg [31:0] dark_weights_normed_update_0_stage_176;
  reg [31:0] dark_weights_normed_update_0_stage_177;
  reg [31:0] dark_weights_normed_update_0_stage_178;
  reg [31:0] dark_weights_normed_update_0_stage_179;
  reg [31:0] dark_weights_normed_update_0_stage_180;
  reg [31:0] dark_weights_normed_update_0_stage_181;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_39;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_40;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_41;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_42;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_43;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_44;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_45;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_46;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_47;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_48;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_49;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_50;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_51;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_52;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_53;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_54;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_55;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_56;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_57;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_58;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_59;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_60;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_61;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_62;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_63;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_64;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_65;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_66;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_67;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_68;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_69;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_70;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_71;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_72;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_73;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_74;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_75;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_76;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_77;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_78;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_79;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_80;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_81;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_82;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_83;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_84;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_85;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_86;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_87;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_88;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_89;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_90;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_91;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_92;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_93;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_94;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_95;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_96;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_97;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_98;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_99;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_100;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_101;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_102;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_103;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_104;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_105;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_106;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_107;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_108;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_109;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_110;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_111;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_112;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_113;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_114;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_115;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_116;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_117;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_118;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_119;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_120;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_121;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_122;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_123;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_124;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_125;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_126;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_127;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_128;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_129;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_130;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_131;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_132;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_133;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_134;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_135;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_136;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_137;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_138;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_139;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_140;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_141;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_142;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_143;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_144;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_145;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_146;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_147;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_148;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_149;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_150;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_151;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_152;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_153;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_154;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_155;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_156;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_157;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_158;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_159;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_160;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_161;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_162;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_163;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_164;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_165;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_166;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_167;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_168;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_169;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_170;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_171;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_172;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_173;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_174;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_175;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_176;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_177;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_178;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_179;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_180;
  reg [287:0] bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_181;
  reg [31:0] bright_gauss_blur_2_update_0_stage_40;
  reg [31:0] bright_gauss_blur_2_update_0_stage_41;
  reg [31:0] bright_gauss_blur_2_update_0_stage_42;
  reg [31:0] bright_gauss_blur_2_update_0_stage_43;
  reg [31:0] bright_gauss_blur_2_update_0_stage_44;
  reg [31:0] bright_gauss_blur_2_update_0_stage_45;
  reg [31:0] bright_gauss_blur_2_update_0_stage_46;
  reg [31:0] bright_gauss_blur_2_update_0_stage_47;
  reg [31:0] bright_gauss_blur_2_update_0_stage_48;
  reg [31:0] bright_gauss_blur_2_update_0_stage_49;
  reg [31:0] bright_gauss_blur_2_update_0_stage_50;
  reg [31:0] bright_gauss_blur_2_update_0_stage_51;
  reg [31:0] bright_gauss_blur_2_update_0_stage_52;
  reg [31:0] bright_gauss_blur_2_update_0_stage_53;
  reg [31:0] bright_gauss_blur_2_update_0_stage_54;
  reg [31:0] bright_gauss_blur_2_update_0_stage_55;
  reg [31:0] bright_gauss_blur_2_update_0_stage_56;
  reg [31:0] bright_gauss_blur_2_update_0_stage_57;
  reg [31:0] bright_gauss_blur_2_update_0_stage_58;
  reg [31:0] bright_gauss_blur_2_update_0_stage_59;
  reg [31:0] bright_gauss_blur_2_update_0_stage_60;
  reg [31:0] bright_gauss_blur_2_update_0_stage_61;
  reg [31:0] bright_gauss_blur_2_update_0_stage_62;
  reg [31:0] bright_gauss_blur_2_update_0_stage_63;
  reg [31:0] bright_gauss_blur_2_update_0_stage_64;
  reg [31:0] bright_gauss_blur_2_update_0_stage_65;
  reg [31:0] bright_gauss_blur_2_update_0_stage_66;
  reg [31:0] bright_gauss_blur_2_update_0_stage_67;
  reg [31:0] bright_gauss_blur_2_update_0_stage_68;
  reg [31:0] bright_gauss_blur_2_update_0_stage_69;
  reg [31:0] bright_gauss_blur_2_update_0_stage_70;
  reg [31:0] bright_gauss_blur_2_update_0_stage_71;
  reg [31:0] bright_gauss_blur_2_update_0_stage_72;
  reg [31:0] bright_gauss_blur_2_update_0_stage_73;
  reg [31:0] bright_gauss_blur_2_update_0_stage_74;
  reg [31:0] bright_gauss_blur_2_update_0_stage_75;
  reg [31:0] bright_gauss_blur_2_update_0_stage_76;
  reg [31:0] bright_gauss_blur_2_update_0_stage_77;
  reg [31:0] bright_gauss_blur_2_update_0_stage_78;
  reg [31:0] bright_gauss_blur_2_update_0_stage_79;
  reg [31:0] bright_gauss_blur_2_update_0_stage_80;
  reg [31:0] bright_gauss_blur_2_update_0_stage_81;
  reg [31:0] bright_gauss_blur_2_update_0_stage_82;
  reg [31:0] bright_gauss_blur_2_update_0_stage_83;
  reg [31:0] bright_gauss_blur_2_update_0_stage_84;
  reg [31:0] bright_gauss_blur_2_update_0_stage_85;
  reg [31:0] bright_gauss_blur_2_update_0_stage_86;
  reg [31:0] bright_gauss_blur_2_update_0_stage_87;
  reg [31:0] bright_gauss_blur_2_update_0_stage_88;
  reg [31:0] bright_gauss_blur_2_update_0_stage_89;
  reg [31:0] bright_gauss_blur_2_update_0_stage_90;
  reg [31:0] bright_gauss_blur_2_update_0_stage_91;
  reg [31:0] bright_gauss_blur_2_update_0_stage_92;
  reg [31:0] bright_gauss_blur_2_update_0_stage_93;
  reg [31:0] bright_gauss_blur_2_update_0_stage_94;
  reg [31:0] bright_gauss_blur_2_update_0_stage_95;
  reg [31:0] bright_gauss_blur_2_update_0_stage_96;
  reg [31:0] bright_gauss_blur_2_update_0_stage_97;
  reg [31:0] bright_gauss_blur_2_update_0_stage_98;
  reg [31:0] bright_gauss_blur_2_update_0_stage_99;
  reg [31:0] bright_gauss_blur_2_update_0_stage_100;
  reg [31:0] bright_gauss_blur_2_update_0_stage_101;
  reg [31:0] bright_gauss_blur_2_update_0_stage_102;
  reg [31:0] bright_gauss_blur_2_update_0_stage_103;
  reg [31:0] bright_gauss_blur_2_update_0_stage_104;
  reg [31:0] bright_gauss_blur_2_update_0_stage_105;
  reg [31:0] bright_gauss_blur_2_update_0_stage_106;
  reg [31:0] bright_gauss_blur_2_update_0_stage_107;
  reg [31:0] bright_gauss_blur_2_update_0_stage_108;
  reg [31:0] bright_gauss_blur_2_update_0_stage_109;
  reg [31:0] bright_gauss_blur_2_update_0_stage_110;
  reg [31:0] bright_gauss_blur_2_update_0_stage_111;
  reg [31:0] bright_gauss_blur_2_update_0_stage_112;
  reg [31:0] bright_gauss_blur_2_update_0_stage_113;
  reg [31:0] bright_gauss_blur_2_update_0_stage_114;
  reg [31:0] bright_gauss_blur_2_update_0_stage_115;
  reg [31:0] bright_gauss_blur_2_update_0_stage_116;
  reg [31:0] bright_gauss_blur_2_update_0_stage_117;
  reg [31:0] bright_gauss_blur_2_update_0_stage_118;
  reg [31:0] bright_gauss_blur_2_update_0_stage_119;
  reg [31:0] bright_gauss_blur_2_update_0_stage_120;
  reg [31:0] bright_gauss_blur_2_update_0_stage_121;
  reg [31:0] bright_gauss_blur_2_update_0_stage_122;
  reg [31:0] bright_gauss_blur_2_update_0_stage_123;
  reg [31:0] bright_gauss_blur_2_update_0_stage_124;
  reg [31:0] bright_gauss_blur_2_update_0_stage_125;
  reg [31:0] bright_gauss_blur_2_update_0_stage_126;
  reg [31:0] bright_gauss_blur_2_update_0_stage_127;
  reg [31:0] bright_gauss_blur_2_update_0_stage_128;
  reg [31:0] bright_gauss_blur_2_update_0_stage_129;
  reg [31:0] bright_gauss_blur_2_update_0_stage_130;
  reg [31:0] bright_gauss_blur_2_update_0_stage_131;
  reg [31:0] bright_gauss_blur_2_update_0_stage_132;
  reg [31:0] bright_gauss_blur_2_update_0_stage_133;
  reg [31:0] bright_gauss_blur_2_update_0_stage_134;
  reg [31:0] bright_gauss_blur_2_update_0_stage_135;
  reg [31:0] bright_gauss_blur_2_update_0_stage_136;
  reg [31:0] bright_gauss_blur_2_update_0_stage_137;
  reg [31:0] bright_gauss_blur_2_update_0_stage_138;
  reg [31:0] bright_gauss_blur_2_update_0_stage_139;
  reg [31:0] bright_gauss_blur_2_update_0_stage_140;
  reg [31:0] bright_gauss_blur_2_update_0_stage_141;
  reg [31:0] bright_gauss_blur_2_update_0_stage_142;
  reg [31:0] bright_gauss_blur_2_update_0_stage_143;
  reg [31:0] bright_gauss_blur_2_update_0_stage_144;
  reg [31:0] bright_gauss_blur_2_update_0_stage_145;
  reg [31:0] bright_gauss_blur_2_update_0_stage_146;
  reg [31:0] bright_gauss_blur_2_update_0_stage_147;
  reg [31:0] bright_gauss_blur_2_update_0_stage_148;
  reg [31:0] bright_gauss_blur_2_update_0_stage_149;
  reg [31:0] bright_gauss_blur_2_update_0_stage_150;
  reg [31:0] bright_gauss_blur_2_update_0_stage_151;
  reg [31:0] bright_gauss_blur_2_update_0_stage_152;
  reg [31:0] bright_gauss_blur_2_update_0_stage_153;
  reg [31:0] bright_gauss_blur_2_update_0_stage_154;
  reg [31:0] bright_gauss_blur_2_update_0_stage_155;
  reg [31:0] bright_gauss_blur_2_update_0_stage_156;
  reg [31:0] bright_gauss_blur_2_update_0_stage_157;
  reg [31:0] bright_gauss_blur_2_update_0_stage_158;
  reg [31:0] bright_gauss_blur_2_update_0_stage_159;
  reg [31:0] bright_gauss_blur_2_update_0_stage_160;
  reg [31:0] bright_gauss_blur_2_update_0_stage_161;
  reg [31:0] bright_gauss_blur_2_update_0_stage_162;
  reg [31:0] bright_gauss_blur_2_update_0_stage_163;
  reg [31:0] bright_gauss_blur_2_update_0_stage_164;
  reg [31:0] bright_gauss_blur_2_update_0_stage_165;
  reg [31:0] bright_gauss_blur_2_update_0_stage_166;
  reg [31:0] bright_gauss_blur_2_update_0_stage_167;
  reg [31:0] bright_gauss_blur_2_update_0_stage_168;
  reg [31:0] bright_gauss_blur_2_update_0_stage_169;
  reg [31:0] bright_gauss_blur_2_update_0_stage_170;
  reg [31:0] bright_gauss_blur_2_update_0_stage_171;
  reg [31:0] bright_gauss_blur_2_update_0_stage_172;
  reg [31:0] bright_gauss_blur_2_update_0_stage_173;
  reg [31:0] bright_gauss_blur_2_update_0_stage_174;
  reg [31:0] bright_gauss_blur_2_update_0_stage_175;
  reg [31:0] bright_gauss_blur_2_update_0_stage_176;
  reg [31:0] bright_gauss_blur_2_update_0_stage_177;
  reg [31:0] bright_gauss_blur_2_update_0_stage_178;
  reg [31:0] bright_gauss_blur_2_update_0_stage_179;
  reg [31:0] bright_gauss_blur_2_update_0_stage_180;
  reg [31:0] bright_gauss_blur_2_update_0_stage_181;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_41;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_42;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_43;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_44;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_45;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_46;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_47;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_48;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_49;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_50;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_51;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_52;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_53;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_54;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_55;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_56;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_57;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_58;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_59;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_60;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_61;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_62;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_63;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_64;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_65;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_66;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_67;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_68;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_69;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_70;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_71;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_72;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_73;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_74;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_75;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_76;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_77;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_78;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_79;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_80;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_81;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_82;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_83;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_84;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_85;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_86;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_87;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_88;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_89;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_90;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_91;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_92;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_93;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_94;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_95;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_96;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_97;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_98;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_99;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_100;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_101;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_102;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_103;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_104;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_105;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_106;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_107;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_108;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_109;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_110;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_111;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_112;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_113;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_114;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_115;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_116;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_117;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_118;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_119;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_120;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_121;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_122;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_123;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_124;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_125;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_126;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_127;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_128;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_129;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_130;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_131;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_132;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_133;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_134;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_135;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_136;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_137;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_138;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_139;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_140;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_141;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_142;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_143;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_144;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_145;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_146;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_147;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_148;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_149;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_150;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_151;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_152;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_153;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_154;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_155;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_156;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_157;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_158;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_159;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_160;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_161;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_162;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_163;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_164;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_165;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_166;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_167;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_168;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_169;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_170;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_171;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_172;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_173;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_174;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_175;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_176;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_177;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_178;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_179;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_180;
  reg [31:0] bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_181;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_46;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_47;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_48;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_49;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_50;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_51;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_52;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_53;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_54;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_55;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_56;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_57;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_58;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_59;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_60;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_61;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_62;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_63;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_64;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_65;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_66;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_67;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_68;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_69;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_70;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_71;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_72;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_73;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_74;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_75;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_76;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_77;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_78;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_79;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_80;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_81;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_82;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_83;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_84;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_85;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_86;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_87;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_88;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_89;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_90;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_91;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_92;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_93;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_94;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_95;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_96;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_97;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_98;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_99;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_100;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_101;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_102;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_103;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_104;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_105;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_106;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_107;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_108;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_109;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_110;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_111;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_112;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_113;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_114;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_115;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_116;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_117;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_118;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_119;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_120;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_121;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_122;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_123;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_124;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_125;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_126;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_127;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_128;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_129;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_130;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_131;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_132;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_133;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_134;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_135;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_136;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_137;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_138;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_139;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_140;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_141;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_142;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_143;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_144;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_145;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_146;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_147;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_148;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_149;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_150;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_151;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_152;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_153;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_154;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_155;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_156;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_157;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_158;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_159;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_160;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_161;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_162;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_163;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_164;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_165;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_166;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_167;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_168;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_169;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_170;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_171;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_172;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_173;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_174;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_175;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_176;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_177;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_178;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_179;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_180;
  reg [31:0] bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_181;
  reg [31:0] bright_laplace_us_0_update_0_stage_47;
  reg [31:0] bright_laplace_us_0_update_0_stage_48;
  reg [31:0] bright_laplace_us_0_update_0_stage_49;
  reg [31:0] bright_laplace_us_0_update_0_stage_50;
  reg [31:0] bright_laplace_us_0_update_0_stage_51;
  reg [31:0] bright_laplace_us_0_update_0_stage_52;
  reg [31:0] bright_laplace_us_0_update_0_stage_53;
  reg [31:0] bright_laplace_us_0_update_0_stage_54;
  reg [31:0] bright_laplace_us_0_update_0_stage_55;
  reg [31:0] bright_laplace_us_0_update_0_stage_56;
  reg [31:0] bright_laplace_us_0_update_0_stage_57;
  reg [31:0] bright_laplace_us_0_update_0_stage_58;
  reg [31:0] bright_laplace_us_0_update_0_stage_59;
  reg [31:0] bright_laplace_us_0_update_0_stage_60;
  reg [31:0] bright_laplace_us_0_update_0_stage_61;
  reg [31:0] bright_laplace_us_0_update_0_stage_62;
  reg [31:0] bright_laplace_us_0_update_0_stage_63;
  reg [31:0] bright_laplace_us_0_update_0_stage_64;
  reg [31:0] bright_laplace_us_0_update_0_stage_65;
  reg [31:0] bright_laplace_us_0_update_0_stage_66;
  reg [31:0] bright_laplace_us_0_update_0_stage_67;
  reg [31:0] bright_laplace_us_0_update_0_stage_68;
  reg [31:0] bright_laplace_us_0_update_0_stage_69;
  reg [31:0] bright_laplace_us_0_update_0_stage_70;
  reg [31:0] bright_laplace_us_0_update_0_stage_71;
  reg [31:0] bright_laplace_us_0_update_0_stage_72;
  reg [31:0] bright_laplace_us_0_update_0_stage_73;
  reg [31:0] bright_laplace_us_0_update_0_stage_74;
  reg [31:0] bright_laplace_us_0_update_0_stage_75;
  reg [31:0] bright_laplace_us_0_update_0_stage_76;
  reg [31:0] bright_laplace_us_0_update_0_stage_77;
  reg [31:0] bright_laplace_us_0_update_0_stage_78;
  reg [31:0] bright_laplace_us_0_update_0_stage_79;
  reg [31:0] bright_laplace_us_0_update_0_stage_80;
  reg [31:0] bright_laplace_us_0_update_0_stage_81;
  reg [31:0] bright_laplace_us_0_update_0_stage_82;
  reg [31:0] bright_laplace_us_0_update_0_stage_83;
  reg [31:0] bright_laplace_us_0_update_0_stage_84;
  reg [31:0] bright_laplace_us_0_update_0_stage_85;
  reg [31:0] bright_laplace_us_0_update_0_stage_86;
  reg [31:0] bright_laplace_us_0_update_0_stage_87;
  reg [31:0] bright_laplace_us_0_update_0_stage_88;
  reg [31:0] bright_laplace_us_0_update_0_stage_89;
  reg [31:0] bright_laplace_us_0_update_0_stage_90;
  reg [31:0] bright_laplace_us_0_update_0_stage_91;
  reg [31:0] bright_laplace_us_0_update_0_stage_92;
  reg [31:0] bright_laplace_us_0_update_0_stage_93;
  reg [31:0] bright_laplace_us_0_update_0_stage_94;
  reg [31:0] bright_laplace_us_0_update_0_stage_95;
  reg [31:0] bright_laplace_us_0_update_0_stage_96;
  reg [31:0] bright_laplace_us_0_update_0_stage_97;
  reg [31:0] bright_laplace_us_0_update_0_stage_98;
  reg [31:0] bright_laplace_us_0_update_0_stage_99;
  reg [31:0] bright_laplace_us_0_update_0_stage_100;
  reg [31:0] bright_laplace_us_0_update_0_stage_101;
  reg [31:0] bright_laplace_us_0_update_0_stage_102;
  reg [31:0] bright_laplace_us_0_update_0_stage_103;
  reg [31:0] bright_laplace_us_0_update_0_stage_104;
  reg [31:0] bright_laplace_us_0_update_0_stage_105;
  reg [31:0] bright_laplace_us_0_update_0_stage_106;
  reg [31:0] bright_laplace_us_0_update_0_stage_107;
  reg [31:0] bright_laplace_us_0_update_0_stage_108;
  reg [31:0] bright_laplace_us_0_update_0_stage_109;
  reg [31:0] bright_laplace_us_0_update_0_stage_110;
  reg [31:0] bright_laplace_us_0_update_0_stage_111;
  reg [31:0] bright_laplace_us_0_update_0_stage_112;
  reg [31:0] bright_laplace_us_0_update_0_stage_113;
  reg [31:0] bright_laplace_us_0_update_0_stage_114;
  reg [31:0] bright_laplace_us_0_update_0_stage_115;
  reg [31:0] bright_laplace_us_0_update_0_stage_116;
  reg [31:0] bright_laplace_us_0_update_0_stage_117;
  reg [31:0] bright_laplace_us_0_update_0_stage_118;
  reg [31:0] bright_laplace_us_0_update_0_stage_119;
  reg [31:0] bright_laplace_us_0_update_0_stage_120;
  reg [31:0] bright_laplace_us_0_update_0_stage_121;
  reg [31:0] bright_laplace_us_0_update_0_stage_122;
  reg [31:0] bright_laplace_us_0_update_0_stage_123;
  reg [31:0] bright_laplace_us_0_update_0_stage_124;
  reg [31:0] bright_laplace_us_0_update_0_stage_125;
  reg [31:0] bright_laplace_us_0_update_0_stage_126;
  reg [31:0] bright_laplace_us_0_update_0_stage_127;
  reg [31:0] bright_laplace_us_0_update_0_stage_128;
  reg [31:0] bright_laplace_us_0_update_0_stage_129;
  reg [31:0] bright_laplace_us_0_update_0_stage_130;
  reg [31:0] bright_laplace_us_0_update_0_stage_131;
  reg [31:0] bright_laplace_us_0_update_0_stage_132;
  reg [31:0] bright_laplace_us_0_update_0_stage_133;
  reg [31:0] bright_laplace_us_0_update_0_stage_134;
  reg [31:0] bright_laplace_us_0_update_0_stage_135;
  reg [31:0] bright_laplace_us_0_update_0_stage_136;
  reg [31:0] bright_laplace_us_0_update_0_stage_137;
  reg [31:0] bright_laplace_us_0_update_0_stage_138;
  reg [31:0] bright_laplace_us_0_update_0_stage_139;
  reg [31:0] bright_laplace_us_0_update_0_stage_140;
  reg [31:0] bright_laplace_us_0_update_0_stage_141;
  reg [31:0] bright_laplace_us_0_update_0_stage_142;
  reg [31:0] bright_laplace_us_0_update_0_stage_143;
  reg [31:0] bright_laplace_us_0_update_0_stage_144;
  reg [31:0] bright_laplace_us_0_update_0_stage_145;
  reg [31:0] bright_laplace_us_0_update_0_stage_146;
  reg [31:0] bright_laplace_us_0_update_0_stage_147;
  reg [31:0] bright_laplace_us_0_update_0_stage_148;
  reg [31:0] bright_laplace_us_0_update_0_stage_149;
  reg [31:0] bright_laplace_us_0_update_0_stage_150;
  reg [31:0] bright_laplace_us_0_update_0_stage_151;
  reg [31:0] bright_laplace_us_0_update_0_stage_152;
  reg [31:0] bright_laplace_us_0_update_0_stage_153;
  reg [31:0] bright_laplace_us_0_update_0_stage_154;
  reg [31:0] bright_laplace_us_0_update_0_stage_155;
  reg [31:0] bright_laplace_us_0_update_0_stage_156;
  reg [31:0] bright_laplace_us_0_update_0_stage_157;
  reg [31:0] bright_laplace_us_0_update_0_stage_158;
  reg [31:0] bright_laplace_us_0_update_0_stage_159;
  reg [31:0] bright_laplace_us_0_update_0_stage_160;
  reg [31:0] bright_laplace_us_0_update_0_stage_161;
  reg [31:0] bright_laplace_us_0_update_0_stage_162;
  reg [31:0] bright_laplace_us_0_update_0_stage_163;
  reg [31:0] bright_laplace_us_0_update_0_stage_164;
  reg [31:0] bright_laplace_us_0_update_0_stage_165;
  reg [31:0] bright_laplace_us_0_update_0_stage_166;
  reg [31:0] bright_laplace_us_0_update_0_stage_167;
  reg [31:0] bright_laplace_us_0_update_0_stage_168;
  reg [31:0] bright_laplace_us_0_update_0_stage_169;
  reg [31:0] bright_laplace_us_0_update_0_stage_170;
  reg [31:0] bright_laplace_us_0_update_0_stage_171;
  reg [31:0] bright_laplace_us_0_update_0_stage_172;
  reg [31:0] bright_laplace_us_0_update_0_stage_173;
  reg [31:0] bright_laplace_us_0_update_0_stage_174;
  reg [31:0] bright_laplace_us_0_update_0_stage_175;
  reg [31:0] bright_laplace_us_0_update_0_stage_176;
  reg [31:0] bright_laplace_us_0_update_0_stage_177;
  reg [31:0] bright_laplace_us_0_update_0_stage_178;
  reg [31:0] bright_laplace_us_0_update_0_stage_179;
  reg [31:0] bright_laplace_us_0_update_0_stage_180;
  reg [31:0] bright_laplace_us_0_update_0_stage_181;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_48;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_49;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_50;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_51;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_52;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_53;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_54;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_55;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_56;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_57;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_58;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_59;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_60;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_61;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_62;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_63;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_64;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_65;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_66;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_67;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_68;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_69;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_70;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_71;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_72;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_73;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_74;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_75;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_76;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_77;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_78;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_79;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_80;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_81;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_82;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_83;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_84;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_85;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_86;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_87;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_88;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_89;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_90;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_91;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_92;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_93;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_94;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_95;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_96;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_97;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_98;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_99;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_100;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_101;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_102;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_103;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_104;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_105;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_106;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_107;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_108;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_109;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_110;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_111;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_112;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_113;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_114;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_115;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_116;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_117;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_118;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_119;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_120;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_121;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_122;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_123;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_124;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_125;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_126;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_127;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_128;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_129;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_130;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_131;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_132;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_133;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_134;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_135;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_136;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_137;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_138;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_139;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_140;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_141;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_142;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_143;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_144;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_145;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_146;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_147;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_148;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_149;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_150;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_151;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_152;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_153;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_154;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_155;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_156;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_157;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_158;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_159;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_160;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_161;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_162;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_163;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_164;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_165;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_166;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_167;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_168;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_169;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_170;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_171;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_172;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_173;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_174;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_175;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_176;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_177;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_178;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_179;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_180;
  reg [31:0] bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_181;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_52;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_53;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_54;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_55;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_56;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_57;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_58;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_59;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_60;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_61;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_62;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_63;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_64;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_65;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_66;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_67;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_68;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_69;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_70;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_71;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_72;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_73;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_74;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_75;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_76;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_77;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_78;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_79;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_80;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_81;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_82;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_83;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_84;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_85;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_86;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_87;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_88;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_89;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_90;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_91;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_92;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_93;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_94;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_95;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_96;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_97;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_98;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_99;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_100;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_101;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_102;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_103;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_104;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_105;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_106;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_107;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_108;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_109;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_110;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_111;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_112;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_113;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_114;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_115;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_116;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_117;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_118;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_119;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_120;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_121;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_122;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_123;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_124;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_125;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_126;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_127;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_128;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_129;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_130;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_131;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_132;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_133;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_134;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_135;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_136;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_137;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_138;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_139;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_140;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_141;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_142;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_143;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_144;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_145;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_146;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_147;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_148;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_149;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_150;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_151;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_152;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_153;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_154;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_155;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_156;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_157;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_158;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_159;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_160;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_161;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_162;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_163;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_164;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_165;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_166;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_167;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_168;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_169;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_170;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_171;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_172;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_173;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_174;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_175;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_176;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_177;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_178;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_179;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_180;
  reg [31:0] dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_181;
  reg [31:0] dark_gauss_ds_2_update_0_stage_53;
  reg [31:0] dark_gauss_ds_2_update_0_stage_54;
  reg [31:0] dark_gauss_ds_2_update_0_stage_55;
  reg [31:0] dark_gauss_ds_2_update_0_stage_56;
  reg [31:0] dark_gauss_ds_2_update_0_stage_57;
  reg [31:0] dark_gauss_ds_2_update_0_stage_58;
  reg [31:0] dark_gauss_ds_2_update_0_stage_59;
  reg [31:0] dark_gauss_ds_2_update_0_stage_60;
  reg [31:0] dark_gauss_ds_2_update_0_stage_61;
  reg [31:0] dark_gauss_ds_2_update_0_stage_62;
  reg [31:0] dark_gauss_ds_2_update_0_stage_63;
  reg [31:0] dark_gauss_ds_2_update_0_stage_64;
  reg [31:0] dark_gauss_ds_2_update_0_stage_65;
  reg [31:0] dark_gauss_ds_2_update_0_stage_66;
  reg [31:0] dark_gauss_ds_2_update_0_stage_67;
  reg [31:0] dark_gauss_ds_2_update_0_stage_68;
  reg [31:0] dark_gauss_ds_2_update_0_stage_69;
  reg [31:0] dark_gauss_ds_2_update_0_stage_70;
  reg [31:0] dark_gauss_ds_2_update_0_stage_71;
  reg [31:0] dark_gauss_ds_2_update_0_stage_72;
  reg [31:0] dark_gauss_ds_2_update_0_stage_73;
  reg [31:0] dark_gauss_ds_2_update_0_stage_74;
  reg [31:0] dark_gauss_ds_2_update_0_stage_75;
  reg [31:0] dark_gauss_ds_2_update_0_stage_76;
  reg [31:0] dark_gauss_ds_2_update_0_stage_77;
  reg [31:0] dark_gauss_ds_2_update_0_stage_78;
  reg [31:0] dark_gauss_ds_2_update_0_stage_79;
  reg [31:0] dark_gauss_ds_2_update_0_stage_80;
  reg [31:0] dark_gauss_ds_2_update_0_stage_81;
  reg [31:0] dark_gauss_ds_2_update_0_stage_82;
  reg [31:0] dark_gauss_ds_2_update_0_stage_83;
  reg [31:0] dark_gauss_ds_2_update_0_stage_84;
  reg [31:0] dark_gauss_ds_2_update_0_stage_85;
  reg [31:0] dark_gauss_ds_2_update_0_stage_86;
  reg [31:0] dark_gauss_ds_2_update_0_stage_87;
  reg [31:0] dark_gauss_ds_2_update_0_stage_88;
  reg [31:0] dark_gauss_ds_2_update_0_stage_89;
  reg [31:0] dark_gauss_ds_2_update_0_stage_90;
  reg [31:0] dark_gauss_ds_2_update_0_stage_91;
  reg [31:0] dark_gauss_ds_2_update_0_stage_92;
  reg [31:0] dark_gauss_ds_2_update_0_stage_93;
  reg [31:0] dark_gauss_ds_2_update_0_stage_94;
  reg [31:0] dark_gauss_ds_2_update_0_stage_95;
  reg [31:0] dark_gauss_ds_2_update_0_stage_96;
  reg [31:0] dark_gauss_ds_2_update_0_stage_97;
  reg [31:0] dark_gauss_ds_2_update_0_stage_98;
  reg [31:0] dark_gauss_ds_2_update_0_stage_99;
  reg [31:0] dark_gauss_ds_2_update_0_stage_100;
  reg [31:0] dark_gauss_ds_2_update_0_stage_101;
  reg [31:0] dark_gauss_ds_2_update_0_stage_102;
  reg [31:0] dark_gauss_ds_2_update_0_stage_103;
  reg [31:0] dark_gauss_ds_2_update_0_stage_104;
  reg [31:0] dark_gauss_ds_2_update_0_stage_105;
  reg [31:0] dark_gauss_ds_2_update_0_stage_106;
  reg [31:0] dark_gauss_ds_2_update_0_stage_107;
  reg [31:0] dark_gauss_ds_2_update_0_stage_108;
  reg [31:0] dark_gauss_ds_2_update_0_stage_109;
  reg [31:0] dark_gauss_ds_2_update_0_stage_110;
  reg [31:0] dark_gauss_ds_2_update_0_stage_111;
  reg [31:0] dark_gauss_ds_2_update_0_stage_112;
  reg [31:0] dark_gauss_ds_2_update_0_stage_113;
  reg [31:0] dark_gauss_ds_2_update_0_stage_114;
  reg [31:0] dark_gauss_ds_2_update_0_stage_115;
  reg [31:0] dark_gauss_ds_2_update_0_stage_116;
  reg [31:0] dark_gauss_ds_2_update_0_stage_117;
  reg [31:0] dark_gauss_ds_2_update_0_stage_118;
  reg [31:0] dark_gauss_ds_2_update_0_stage_119;
  reg [31:0] dark_gauss_ds_2_update_0_stage_120;
  reg [31:0] dark_gauss_ds_2_update_0_stage_121;
  reg [31:0] dark_gauss_ds_2_update_0_stage_122;
  reg [31:0] dark_gauss_ds_2_update_0_stage_123;
  reg [31:0] dark_gauss_ds_2_update_0_stage_124;
  reg [31:0] dark_gauss_ds_2_update_0_stage_125;
  reg [31:0] dark_gauss_ds_2_update_0_stage_126;
  reg [31:0] dark_gauss_ds_2_update_0_stage_127;
  reg [31:0] dark_gauss_ds_2_update_0_stage_128;
  reg [31:0] dark_gauss_ds_2_update_0_stage_129;
  reg [31:0] dark_gauss_ds_2_update_0_stage_130;
  reg [31:0] dark_gauss_ds_2_update_0_stage_131;
  reg [31:0] dark_gauss_ds_2_update_0_stage_132;
  reg [31:0] dark_gauss_ds_2_update_0_stage_133;
  reg [31:0] dark_gauss_ds_2_update_0_stage_134;
  reg [31:0] dark_gauss_ds_2_update_0_stage_135;
  reg [31:0] dark_gauss_ds_2_update_0_stage_136;
  reg [31:0] dark_gauss_ds_2_update_0_stage_137;
  reg [31:0] dark_gauss_ds_2_update_0_stage_138;
  reg [31:0] dark_gauss_ds_2_update_0_stage_139;
  reg [31:0] dark_gauss_ds_2_update_0_stage_140;
  reg [31:0] dark_gauss_ds_2_update_0_stage_141;
  reg [31:0] dark_gauss_ds_2_update_0_stage_142;
  reg [31:0] dark_gauss_ds_2_update_0_stage_143;
  reg [31:0] dark_gauss_ds_2_update_0_stage_144;
  reg [31:0] dark_gauss_ds_2_update_0_stage_145;
  reg [31:0] dark_gauss_ds_2_update_0_stage_146;
  reg [31:0] dark_gauss_ds_2_update_0_stage_147;
  reg [31:0] dark_gauss_ds_2_update_0_stage_148;
  reg [31:0] dark_gauss_ds_2_update_0_stage_149;
  reg [31:0] dark_gauss_ds_2_update_0_stage_150;
  reg [31:0] dark_gauss_ds_2_update_0_stage_151;
  reg [31:0] dark_gauss_ds_2_update_0_stage_152;
  reg [31:0] dark_gauss_ds_2_update_0_stage_153;
  reg [31:0] dark_gauss_ds_2_update_0_stage_154;
  reg [31:0] dark_gauss_ds_2_update_0_stage_155;
  reg [31:0] dark_gauss_ds_2_update_0_stage_156;
  reg [31:0] dark_gauss_ds_2_update_0_stage_157;
  reg [31:0] dark_gauss_ds_2_update_0_stage_158;
  reg [31:0] dark_gauss_ds_2_update_0_stage_159;
  reg [31:0] dark_gauss_ds_2_update_0_stage_160;
  reg [31:0] dark_gauss_ds_2_update_0_stage_161;
  reg [31:0] dark_gauss_ds_2_update_0_stage_162;
  reg [31:0] dark_gauss_ds_2_update_0_stage_163;
  reg [31:0] dark_gauss_ds_2_update_0_stage_164;
  reg [31:0] dark_gauss_ds_2_update_0_stage_165;
  reg [31:0] dark_gauss_ds_2_update_0_stage_166;
  reg [31:0] dark_gauss_ds_2_update_0_stage_167;
  reg [31:0] dark_gauss_ds_2_update_0_stage_168;
  reg [31:0] dark_gauss_ds_2_update_0_stage_169;
  reg [31:0] dark_gauss_ds_2_update_0_stage_170;
  reg [31:0] dark_gauss_ds_2_update_0_stage_171;
  reg [31:0] dark_gauss_ds_2_update_0_stage_172;
  reg [31:0] dark_gauss_ds_2_update_0_stage_173;
  reg [31:0] dark_gauss_ds_2_update_0_stage_174;
  reg [31:0] dark_gauss_ds_2_update_0_stage_175;
  reg [31:0] dark_gauss_ds_2_update_0_stage_176;
  reg [31:0] dark_gauss_ds_2_update_0_stage_177;
  reg [31:0] dark_gauss_ds_2_update_0_stage_178;
  reg [31:0] dark_gauss_ds_2_update_0_stage_179;
  reg [31:0] dark_gauss_ds_2_update_0_stage_180;
  reg [31:0] dark_gauss_ds_2_update_0_stage_181;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_54;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_55;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_56;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_57;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_58;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_59;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_60;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_61;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_62;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_63;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_64;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_65;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_66;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_67;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_68;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_69;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_70;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_71;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_72;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_73;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_74;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_75;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_76;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_77;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_78;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_79;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_80;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_81;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_82;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_83;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_84;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_85;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_86;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_87;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_88;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_89;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_90;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_91;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_92;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_93;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_94;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_95;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_96;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_97;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_98;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_99;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_100;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_101;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_102;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_103;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_104;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_105;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_106;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_107;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_108;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_109;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_110;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_111;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_112;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_113;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_114;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_115;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_116;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_117;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_118;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_119;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_120;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_121;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_122;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_123;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_124;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_125;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_126;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_127;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_128;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_129;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_130;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_131;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_132;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_133;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_134;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_135;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_136;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_137;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_138;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_139;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_140;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_141;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_142;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_143;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_144;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_145;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_146;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_147;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_148;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_149;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_150;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_151;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_152;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_153;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_154;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_155;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_156;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_157;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_158;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_159;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_160;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_161;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_162;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_163;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_164;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_165;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_166;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_167;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_168;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_169;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_170;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_171;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_172;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_173;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_174;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_175;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_176;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_177;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_178;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_179;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_180;
  reg [31:0] dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_181;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_107;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_108;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_109;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_110;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_111;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_112;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_113;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_114;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_115;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_116;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_117;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_118;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_119;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_120;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_121;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_122;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_123;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_124;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_125;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_126;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_127;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_128;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_129;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_130;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_131;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_132;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_133;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_134;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_135;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_136;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_137;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_138;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_139;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_140;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_141;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_142;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_143;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_144;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_145;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_146;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_147;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_148;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_149;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_150;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_151;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_152;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_153;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_154;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_155;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_156;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_157;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_158;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_159;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_160;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_161;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_162;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_163;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_164;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_165;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_166;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_167;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_168;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_169;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_170;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_171;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_172;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_173;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_174;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_175;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_176;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_177;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_178;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_179;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_180;
  reg [287:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_181;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_55;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_56;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_57;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_58;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_59;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_60;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_61;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_62;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_63;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_64;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_65;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_66;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_67;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_68;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_69;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_70;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_71;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_72;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_73;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_74;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_75;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_76;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_77;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_78;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_79;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_80;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_81;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_82;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_83;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_84;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_85;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_86;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_87;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_88;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_89;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_90;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_91;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_92;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_93;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_94;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_95;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_96;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_97;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_98;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_99;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_100;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_101;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_102;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_103;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_104;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_105;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_106;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_107;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_108;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_109;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_110;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_111;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_112;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_113;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_114;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_115;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_116;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_117;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_118;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_119;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_120;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_121;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_122;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_123;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_124;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_125;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_126;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_127;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_128;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_129;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_130;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_131;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_132;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_133;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_134;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_135;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_136;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_137;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_138;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_139;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_140;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_141;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_142;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_143;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_144;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_145;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_146;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_147;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_148;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_149;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_150;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_151;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_152;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_153;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_154;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_155;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_156;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_157;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_158;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_159;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_160;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_161;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_162;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_163;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_164;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_165;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_166;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_167;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_168;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_169;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_170;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_171;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_172;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_173;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_174;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_175;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_176;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_177;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_178;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_179;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_180;
  reg [287:0] bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_181;
  reg [31:0] bright_gauss_blur_3_update_0_stage_56;
  reg [31:0] bright_gauss_blur_3_update_0_stage_57;
  reg [31:0] bright_gauss_blur_3_update_0_stage_58;
  reg [31:0] bright_gauss_blur_3_update_0_stage_59;
  reg [31:0] bright_gauss_blur_3_update_0_stage_60;
  reg [31:0] bright_gauss_blur_3_update_0_stage_61;
  reg [31:0] bright_gauss_blur_3_update_0_stage_62;
  reg [31:0] bright_gauss_blur_3_update_0_stage_63;
  reg [31:0] bright_gauss_blur_3_update_0_stage_64;
  reg [31:0] bright_gauss_blur_3_update_0_stage_65;
  reg [31:0] bright_gauss_blur_3_update_0_stage_66;
  reg [31:0] bright_gauss_blur_3_update_0_stage_67;
  reg [31:0] bright_gauss_blur_3_update_0_stage_68;
  reg [31:0] bright_gauss_blur_3_update_0_stage_69;
  reg [31:0] bright_gauss_blur_3_update_0_stage_70;
  reg [31:0] bright_gauss_blur_3_update_0_stage_71;
  reg [31:0] bright_gauss_blur_3_update_0_stage_72;
  reg [31:0] bright_gauss_blur_3_update_0_stage_73;
  reg [31:0] bright_gauss_blur_3_update_0_stage_74;
  reg [31:0] bright_gauss_blur_3_update_0_stage_75;
  reg [31:0] bright_gauss_blur_3_update_0_stage_76;
  reg [31:0] bright_gauss_blur_3_update_0_stage_77;
  reg [31:0] bright_gauss_blur_3_update_0_stage_78;
  reg [31:0] bright_gauss_blur_3_update_0_stage_79;
  reg [31:0] bright_gauss_blur_3_update_0_stage_80;
  reg [31:0] bright_gauss_blur_3_update_0_stage_81;
  reg [31:0] bright_gauss_blur_3_update_0_stage_82;
  reg [31:0] bright_gauss_blur_3_update_0_stage_83;
  reg [31:0] bright_gauss_blur_3_update_0_stage_84;
  reg [31:0] bright_gauss_blur_3_update_0_stage_85;
  reg [31:0] bright_gauss_blur_3_update_0_stage_86;
  reg [31:0] bright_gauss_blur_3_update_0_stage_87;
  reg [31:0] bright_gauss_blur_3_update_0_stage_88;
  reg [31:0] bright_gauss_blur_3_update_0_stage_89;
  reg [31:0] bright_gauss_blur_3_update_0_stage_90;
  reg [31:0] bright_gauss_blur_3_update_0_stage_91;
  reg [31:0] bright_gauss_blur_3_update_0_stage_92;
  reg [31:0] bright_gauss_blur_3_update_0_stage_93;
  reg [31:0] bright_gauss_blur_3_update_0_stage_94;
  reg [31:0] bright_gauss_blur_3_update_0_stage_95;
  reg [31:0] bright_gauss_blur_3_update_0_stage_96;
  reg [31:0] bright_gauss_blur_3_update_0_stage_97;
  reg [31:0] bright_gauss_blur_3_update_0_stage_98;
  reg [31:0] bright_gauss_blur_3_update_0_stage_99;
  reg [31:0] bright_gauss_blur_3_update_0_stage_100;
  reg [31:0] bright_gauss_blur_3_update_0_stage_101;
  reg [31:0] bright_gauss_blur_3_update_0_stage_102;
  reg [31:0] bright_gauss_blur_3_update_0_stage_103;
  reg [31:0] bright_gauss_blur_3_update_0_stage_104;
  reg [31:0] bright_gauss_blur_3_update_0_stage_105;
  reg [31:0] bright_gauss_blur_3_update_0_stage_106;
  reg [31:0] bright_gauss_blur_3_update_0_stage_107;
  reg [31:0] bright_gauss_blur_3_update_0_stage_108;
  reg [31:0] bright_gauss_blur_3_update_0_stage_109;
  reg [31:0] bright_gauss_blur_3_update_0_stage_110;
  reg [31:0] bright_gauss_blur_3_update_0_stage_111;
  reg [31:0] bright_gauss_blur_3_update_0_stage_112;
  reg [31:0] bright_gauss_blur_3_update_0_stage_113;
  reg [31:0] bright_gauss_blur_3_update_0_stage_114;
  reg [31:0] bright_gauss_blur_3_update_0_stage_115;
  reg [31:0] bright_gauss_blur_3_update_0_stage_116;
  reg [31:0] bright_gauss_blur_3_update_0_stage_117;
  reg [31:0] bright_gauss_blur_3_update_0_stage_118;
  reg [31:0] bright_gauss_blur_3_update_0_stage_119;
  reg [31:0] bright_gauss_blur_3_update_0_stage_120;
  reg [31:0] bright_gauss_blur_3_update_0_stage_121;
  reg [31:0] bright_gauss_blur_3_update_0_stage_122;
  reg [31:0] bright_gauss_blur_3_update_0_stage_123;
  reg [31:0] bright_gauss_blur_3_update_0_stage_124;
  reg [31:0] bright_gauss_blur_3_update_0_stage_125;
  reg [31:0] bright_gauss_blur_3_update_0_stage_126;
  reg [31:0] bright_gauss_blur_3_update_0_stage_127;
  reg [31:0] bright_gauss_blur_3_update_0_stage_128;
  reg [31:0] bright_gauss_blur_3_update_0_stage_129;
  reg [31:0] bright_gauss_blur_3_update_0_stage_130;
  reg [31:0] bright_gauss_blur_3_update_0_stage_131;
  reg [31:0] bright_gauss_blur_3_update_0_stage_132;
  reg [31:0] bright_gauss_blur_3_update_0_stage_133;
  reg [31:0] bright_gauss_blur_3_update_0_stage_134;
  reg [31:0] bright_gauss_blur_3_update_0_stage_135;
  reg [31:0] bright_gauss_blur_3_update_0_stage_136;
  reg [31:0] bright_gauss_blur_3_update_0_stage_137;
  reg [31:0] bright_gauss_blur_3_update_0_stage_138;
  reg [31:0] bright_gauss_blur_3_update_0_stage_139;
  reg [31:0] bright_gauss_blur_3_update_0_stage_140;
  reg [31:0] bright_gauss_blur_3_update_0_stage_141;
  reg [31:0] bright_gauss_blur_3_update_0_stage_142;
  reg [31:0] bright_gauss_blur_3_update_0_stage_143;
  reg [31:0] bright_gauss_blur_3_update_0_stage_144;
  reg [31:0] bright_gauss_blur_3_update_0_stage_145;
  reg [31:0] bright_gauss_blur_3_update_0_stage_146;
  reg [31:0] bright_gauss_blur_3_update_0_stage_147;
  reg [31:0] bright_gauss_blur_3_update_0_stage_148;
  reg [31:0] bright_gauss_blur_3_update_0_stage_149;
  reg [31:0] bright_gauss_blur_3_update_0_stage_150;
  reg [31:0] bright_gauss_blur_3_update_0_stage_151;
  reg [31:0] bright_gauss_blur_3_update_0_stage_152;
  reg [31:0] bright_gauss_blur_3_update_0_stage_153;
  reg [31:0] bright_gauss_blur_3_update_0_stage_154;
  reg [31:0] bright_gauss_blur_3_update_0_stage_155;
  reg [31:0] bright_gauss_blur_3_update_0_stage_156;
  reg [31:0] bright_gauss_blur_3_update_0_stage_157;
  reg [31:0] bright_gauss_blur_3_update_0_stage_158;
  reg [31:0] bright_gauss_blur_3_update_0_stage_159;
  reg [31:0] bright_gauss_blur_3_update_0_stage_160;
  reg [31:0] bright_gauss_blur_3_update_0_stage_161;
  reg [31:0] bright_gauss_blur_3_update_0_stage_162;
  reg [31:0] bright_gauss_blur_3_update_0_stage_163;
  reg [31:0] bright_gauss_blur_3_update_0_stage_164;
  reg [31:0] bright_gauss_blur_3_update_0_stage_165;
  reg [31:0] bright_gauss_blur_3_update_0_stage_166;
  reg [31:0] bright_gauss_blur_3_update_0_stage_167;
  reg [31:0] bright_gauss_blur_3_update_0_stage_168;
  reg [31:0] bright_gauss_blur_3_update_0_stage_169;
  reg [31:0] bright_gauss_blur_3_update_0_stage_170;
  reg [31:0] bright_gauss_blur_3_update_0_stage_171;
  reg [31:0] bright_gauss_blur_3_update_0_stage_172;
  reg [31:0] bright_gauss_blur_3_update_0_stage_173;
  reg [31:0] bright_gauss_blur_3_update_0_stage_174;
  reg [31:0] bright_gauss_blur_3_update_0_stage_175;
  reg [31:0] bright_gauss_blur_3_update_0_stage_176;
  reg [31:0] bright_gauss_blur_3_update_0_stage_177;
  reg [31:0] bright_gauss_blur_3_update_0_stage_178;
  reg [31:0] bright_gauss_blur_3_update_0_stage_179;
  reg [31:0] bright_gauss_blur_3_update_0_stage_180;
  reg [31:0] bright_gauss_blur_3_update_0_stage_181;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_57;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_58;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_59;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_60;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_61;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_62;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_63;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_64;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_65;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_66;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_67;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_68;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_69;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_70;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_71;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_72;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_73;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_74;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_75;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_76;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_77;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_78;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_79;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_80;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_81;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_82;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_83;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_84;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_85;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_86;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_87;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_88;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_89;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_90;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_91;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_92;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_93;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_94;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_95;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_96;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_97;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_98;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_99;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_100;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_101;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_102;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_103;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_104;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_105;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_106;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_107;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_108;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_109;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_110;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_111;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_112;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_113;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_114;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_115;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_116;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_117;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_118;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_119;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_120;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_121;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_122;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_123;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_124;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_125;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_126;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_127;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_128;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_129;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_130;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_131;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_132;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_133;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_134;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_135;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_136;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_137;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_138;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_139;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_140;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_141;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_142;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_143;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_144;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_145;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_146;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_147;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_148;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_149;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_150;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_151;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_152;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_153;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_154;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_155;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_156;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_157;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_158;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_159;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_160;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_161;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_162;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_163;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_164;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_165;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_166;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_167;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_168;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_169;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_170;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_171;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_172;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_173;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_174;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_175;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_176;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_177;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_178;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_179;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_180;
  reg [31:0] bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_181;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_68;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_69;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_70;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_71;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_72;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_73;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_74;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_75;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_76;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_77;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_78;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_79;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_80;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_81;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_82;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_83;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_84;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_85;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_86;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_87;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_88;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_89;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_90;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_91;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_92;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_93;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_94;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_95;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_96;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_97;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_98;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_99;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_100;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_101;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_102;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_103;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_104;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_105;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_106;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_107;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_108;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_109;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_110;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_111;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_112;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_113;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_114;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_115;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_116;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_117;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_118;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_119;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_120;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_121;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_122;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_123;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_124;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_125;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_126;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_127;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_128;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_129;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_130;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_131;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_132;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_133;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_134;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_135;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_136;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_137;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_138;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_139;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_140;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_141;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_142;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_143;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_144;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_145;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_146;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_147;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_148;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_149;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_150;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_151;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_152;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_153;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_154;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_155;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_156;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_157;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_158;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_159;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_160;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_161;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_162;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_163;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_164;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_165;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_166;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_167;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_168;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_169;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_170;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_171;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_172;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_173;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_174;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_175;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_176;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_177;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_178;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_179;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_180;
  reg [31:0] dark_weights_dark_weights_normed_update_0_read_read_45_stage_181;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_71;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_72;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_73;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_74;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_75;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_76;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_77;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_78;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_79;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_80;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_81;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_82;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_83;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_84;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_85;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_86;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_87;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_88;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_89;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_90;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_91;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_92;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_93;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_94;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_95;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_96;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_97;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_98;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_99;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_100;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_101;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_102;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_103;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_104;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_105;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_106;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_107;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_108;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_109;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_110;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_111;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_112;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_113;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_114;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_115;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_116;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_117;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_118;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_119;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_120;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_121;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_122;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_123;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_124;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_125;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_126;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_127;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_128;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_129;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_130;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_131;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_132;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_133;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_134;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_135;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_136;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_137;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_138;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_139;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_140;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_141;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_142;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_143;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_144;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_145;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_146;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_147;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_148;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_149;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_150;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_151;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_152;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_153;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_154;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_155;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_156;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_157;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_158;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_159;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_160;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_161;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_162;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_163;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_164;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_165;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_166;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_167;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_168;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_169;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_170;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_171;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_172;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_173;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_174;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_175;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_176;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_177;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_178;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_179;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_180;
  reg [31:0] dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_181;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_76;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_77;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_78;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_79;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_80;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_81;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_82;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_83;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_84;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_85;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_86;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_87;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_88;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_89;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_90;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_91;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_92;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_93;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_94;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_95;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_96;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_97;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_98;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_99;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_100;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_101;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_102;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_103;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_104;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_105;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_106;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_107;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_108;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_109;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_110;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_111;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_112;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_113;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_114;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_115;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_116;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_117;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_118;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_119;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_120;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_121;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_122;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_123;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_124;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_125;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_126;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_127;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_128;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_129;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_130;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_131;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_132;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_133;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_134;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_135;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_136;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_137;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_138;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_139;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_140;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_141;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_142;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_143;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_144;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_145;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_146;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_147;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_148;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_149;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_150;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_151;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_152;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_153;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_154;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_155;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_156;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_157;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_158;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_159;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_160;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_161;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_162;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_163;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_164;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_165;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_166;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_167;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_168;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_169;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_170;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_171;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_172;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_173;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_174;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_175;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_176;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_177;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_178;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_179;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_180;
  reg [287:0] dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_77;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_78;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_79;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_80;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_81;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_82;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_83;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_84;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_85;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_86;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_87;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_88;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_89;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_90;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_91;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_92;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_93;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_1_update_0_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_78;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_79;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_80;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_81;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_82;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_83;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_84;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_85;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_86;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_87;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_88;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_89;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_90;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_91;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_92;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_93;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_181;
  reg [31:0] dark_laplace_us_1_update_0_stage_92;
  reg [31:0] dark_laplace_us_1_update_0_stage_93;
  reg [31:0] dark_laplace_us_1_update_0_stage_94;
  reg [31:0] dark_laplace_us_1_update_0_stage_95;
  reg [31:0] dark_laplace_us_1_update_0_stage_96;
  reg [31:0] dark_laplace_us_1_update_0_stage_97;
  reg [31:0] dark_laplace_us_1_update_0_stage_98;
  reg [31:0] dark_laplace_us_1_update_0_stage_99;
  reg [31:0] dark_laplace_us_1_update_0_stage_100;
  reg [31:0] dark_laplace_us_1_update_0_stage_101;
  reg [31:0] dark_laplace_us_1_update_0_stage_102;
  reg [31:0] dark_laplace_us_1_update_0_stage_103;
  reg [31:0] dark_laplace_us_1_update_0_stage_104;
  reg [31:0] dark_laplace_us_1_update_0_stage_105;
  reg [31:0] dark_laplace_us_1_update_0_stage_106;
  reg [31:0] dark_laplace_us_1_update_0_stage_107;
  reg [31:0] dark_laplace_us_1_update_0_stage_108;
  reg [31:0] dark_laplace_us_1_update_0_stage_109;
  reg [31:0] dark_laplace_us_1_update_0_stage_110;
  reg [31:0] dark_laplace_us_1_update_0_stage_111;
  reg [31:0] dark_laplace_us_1_update_0_stage_112;
  reg [31:0] dark_laplace_us_1_update_0_stage_113;
  reg [31:0] dark_laplace_us_1_update_0_stage_114;
  reg [31:0] dark_laplace_us_1_update_0_stage_115;
  reg [31:0] dark_laplace_us_1_update_0_stage_116;
  reg [31:0] dark_laplace_us_1_update_0_stage_117;
  reg [31:0] dark_laplace_us_1_update_0_stage_118;
  reg [31:0] dark_laplace_us_1_update_0_stage_119;
  reg [31:0] dark_laplace_us_1_update_0_stage_120;
  reg [31:0] dark_laplace_us_1_update_0_stage_121;
  reg [31:0] dark_laplace_us_1_update_0_stage_122;
  reg [31:0] dark_laplace_us_1_update_0_stage_123;
  reg [31:0] dark_laplace_us_1_update_0_stage_124;
  reg [31:0] dark_laplace_us_1_update_0_stage_125;
  reg [31:0] dark_laplace_us_1_update_0_stage_126;
  reg [31:0] dark_laplace_us_1_update_0_stage_127;
  reg [31:0] dark_laplace_us_1_update_0_stage_128;
  reg [31:0] dark_laplace_us_1_update_0_stage_129;
  reg [31:0] dark_laplace_us_1_update_0_stage_130;
  reg [31:0] dark_laplace_us_1_update_0_stage_131;
  reg [31:0] dark_laplace_us_1_update_0_stage_132;
  reg [31:0] dark_laplace_us_1_update_0_stage_133;
  reg [31:0] dark_laplace_us_1_update_0_stage_134;
  reg [31:0] dark_laplace_us_1_update_0_stage_135;
  reg [31:0] dark_laplace_us_1_update_0_stage_136;
  reg [31:0] dark_laplace_us_1_update_0_stage_137;
  reg [31:0] dark_laplace_us_1_update_0_stage_138;
  reg [31:0] dark_laplace_us_1_update_0_stage_139;
  reg [31:0] dark_laplace_us_1_update_0_stage_140;
  reg [31:0] dark_laplace_us_1_update_0_stage_141;
  reg [31:0] dark_laplace_us_1_update_0_stage_142;
  reg [31:0] dark_laplace_us_1_update_0_stage_143;
  reg [31:0] dark_laplace_us_1_update_0_stage_144;
  reg [31:0] dark_laplace_us_1_update_0_stage_145;
  reg [31:0] dark_laplace_us_1_update_0_stage_146;
  reg [31:0] dark_laplace_us_1_update_0_stage_147;
  reg [31:0] dark_laplace_us_1_update_0_stage_148;
  reg [31:0] dark_laplace_us_1_update_0_stage_149;
  reg [31:0] dark_laplace_us_1_update_0_stage_150;
  reg [31:0] dark_laplace_us_1_update_0_stage_151;
  reg [31:0] dark_laplace_us_1_update_0_stage_152;
  reg [31:0] dark_laplace_us_1_update_0_stage_153;
  reg [31:0] dark_laplace_us_1_update_0_stage_154;
  reg [31:0] dark_laplace_us_1_update_0_stage_155;
  reg [31:0] dark_laplace_us_1_update_0_stage_156;
  reg [31:0] dark_laplace_us_1_update_0_stage_157;
  reg [31:0] dark_laplace_us_1_update_0_stage_158;
  reg [31:0] dark_laplace_us_1_update_0_stage_159;
  reg [31:0] dark_laplace_us_1_update_0_stage_160;
  reg [31:0] dark_laplace_us_1_update_0_stage_161;
  reg [31:0] dark_laplace_us_1_update_0_stage_162;
  reg [31:0] dark_laplace_us_1_update_0_stage_163;
  reg [31:0] dark_laplace_us_1_update_0_stage_164;
  reg [31:0] dark_laplace_us_1_update_0_stage_165;
  reg [31:0] dark_laplace_us_1_update_0_stage_166;
  reg [31:0] dark_laplace_us_1_update_0_stage_167;
  reg [31:0] dark_laplace_us_1_update_0_stage_168;
  reg [31:0] dark_laplace_us_1_update_0_stage_169;
  reg [31:0] dark_laplace_us_1_update_0_stage_170;
  reg [31:0] dark_laplace_us_1_update_0_stage_171;
  reg [31:0] dark_laplace_us_1_update_0_stage_172;
  reg [31:0] dark_laplace_us_1_update_0_stage_173;
  reg [31:0] dark_laplace_us_1_update_0_stage_174;
  reg [31:0] dark_laplace_us_1_update_0_stage_175;
  reg [31:0] dark_laplace_us_1_update_0_stage_176;
  reg [31:0] dark_laplace_us_1_update_0_stage_177;
  reg [31:0] dark_laplace_us_1_update_0_stage_178;
  reg [31:0] dark_laplace_us_1_update_0_stage_179;
  reg [31:0] dark_laplace_us_1_update_0_stage_180;
  reg [31:0] dark_laplace_us_1_update_0_stage_181;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_93;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_94;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_95;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_96;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_97;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_98;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_99;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_100;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_101;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_102;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_103;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_104;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_105;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_106;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_107;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_108;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_109;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_110;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_111;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_112;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_113;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_114;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_115;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_116;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_117;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_118;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_119;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_120;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_121;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_122;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_123;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_124;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_125;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_126;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_127;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_128;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_129;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_130;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_131;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_132;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_133;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_134;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_135;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_136;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_137;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_138;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_139;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_140;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_141;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_142;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_143;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_144;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_145;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_146;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_147;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_148;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_149;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_150;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_151;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_152;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_153;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_154;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_155;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_156;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_157;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_158;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_159;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_160;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_161;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_162;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_163;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_164;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_165;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_166;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_167;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_168;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_169;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_170;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_171;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_172;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_173;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_174;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_175;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_176;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_177;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_178;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_179;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_180;
  reg [31:0] dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_181;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_100;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_101;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_102;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_103;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_104;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_105;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_106;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_107;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_108;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_109;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_110;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_111;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_112;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_113;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_114;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_115;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_116;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_117;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_118;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_119;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_120;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_121;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_122;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_123;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_124;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_125;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_126;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_127;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_128;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_129;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_130;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_131;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_132;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_133;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_134;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_135;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_136;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_137;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_138;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_139;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_140;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_141;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_142;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_143;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_144;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_145;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_146;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_147;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_148;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_149;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_150;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_151;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_152;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_153;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_154;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_155;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_156;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_157;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_158;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_159;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_160;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_161;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_162;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_163;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_164;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_165;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_166;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_167;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_168;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_169;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_170;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_171;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_172;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_173;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_174;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_175;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_176;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_177;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_178;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_179;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_180;
  reg [31:0] bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_94;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_95;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_96;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_97;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_98;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_99;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_100;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_101;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_102;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_103;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_104;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_105;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_106;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_107;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_95;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_96;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_97;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_98;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_99;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_100;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_101;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_102;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_103;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_104;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_105;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_106;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_107;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_108;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_109;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_110;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_111;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_112;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_113;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_114;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_115;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_116;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_117;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_118;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_119;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_120;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_121;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_122;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_123;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_124;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_125;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_126;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_127;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_128;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_129;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_130;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_131;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_132;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_133;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_134;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_135;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_136;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_2_update_0_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_96;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_97;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_98;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_99;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_100;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_101;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_102;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_103;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_104;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_105;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_106;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_107;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_108;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_109;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_110;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_111;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_112;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_113;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_114;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_115;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_116;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_117;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_118;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_119;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_120;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_121;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_122;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_123;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_124;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_125;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_126;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_127;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_128;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_129;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_130;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_131;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_132;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_133;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_134;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_135;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_136;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_137;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_138;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_139;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_140;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_141;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_142;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_143;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_144;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_145;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_146;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_147;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_148;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_149;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_150;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_151;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_152;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_153;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_154;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_155;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_156;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_157;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_181;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_101;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_102;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_103;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_104;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_105;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_106;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_107;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_108;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_109;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_110;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_111;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_112;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_113;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_114;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_115;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_116;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_117;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_118;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_119;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_120;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_121;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_122;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_123;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_124;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_125;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_126;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_127;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_128;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_129;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_130;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_131;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_132;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_133;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_134;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_135;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_136;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_137;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_138;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_139;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_140;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_141;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_142;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_143;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_144;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_145;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_146;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_147;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_148;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_149;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_150;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_151;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_152;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_153;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_154;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_155;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_156;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_157;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_158;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_159;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_160;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_161;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_162;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_163;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_164;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_165;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_166;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_167;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_168;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_169;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_170;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_171;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_172;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_173;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_174;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_175;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_176;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_177;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_178;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_179;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_180;
  reg [31:0] bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_181;
  reg [31:0] bright_laplace_diff_1_update_0_stage_102;
  reg [31:0] bright_laplace_diff_1_update_0_stage_103;
  reg [31:0] bright_laplace_diff_1_update_0_stage_104;
  reg [31:0] bright_laplace_diff_1_update_0_stage_105;
  reg [31:0] bright_laplace_diff_1_update_0_stage_106;
  reg [31:0] bright_laplace_diff_1_update_0_stage_107;
  reg [31:0] bright_laplace_diff_1_update_0_stage_108;
  reg [31:0] bright_laplace_diff_1_update_0_stage_109;
  reg [31:0] bright_laplace_diff_1_update_0_stage_110;
  reg [31:0] bright_laplace_diff_1_update_0_stage_111;
  reg [31:0] bright_laplace_diff_1_update_0_stage_112;
  reg [31:0] bright_laplace_diff_1_update_0_stage_113;
  reg [31:0] bright_laplace_diff_1_update_0_stage_114;
  reg [31:0] bright_laplace_diff_1_update_0_stage_115;
  reg [31:0] bright_laplace_diff_1_update_0_stage_116;
  reg [31:0] bright_laplace_diff_1_update_0_stage_117;
  reg [31:0] bright_laplace_diff_1_update_0_stage_118;
  reg [31:0] bright_laplace_diff_1_update_0_stage_119;
  reg [31:0] bright_laplace_diff_1_update_0_stage_120;
  reg [31:0] bright_laplace_diff_1_update_0_stage_121;
  reg [31:0] bright_laplace_diff_1_update_0_stage_122;
  reg [31:0] bright_laplace_diff_1_update_0_stage_123;
  reg [31:0] bright_laplace_diff_1_update_0_stage_124;
  reg [31:0] bright_laplace_diff_1_update_0_stage_125;
  reg [31:0] bright_laplace_diff_1_update_0_stage_126;
  reg [31:0] bright_laplace_diff_1_update_0_stage_127;
  reg [31:0] bright_laplace_diff_1_update_0_stage_128;
  reg [31:0] bright_laplace_diff_1_update_0_stage_129;
  reg [31:0] bright_laplace_diff_1_update_0_stage_130;
  reg [31:0] bright_laplace_diff_1_update_0_stage_131;
  reg [31:0] bright_laplace_diff_1_update_0_stage_132;
  reg [31:0] bright_laplace_diff_1_update_0_stage_133;
  reg [31:0] bright_laplace_diff_1_update_0_stage_134;
  reg [31:0] bright_laplace_diff_1_update_0_stage_135;
  reg [31:0] bright_laplace_diff_1_update_0_stage_136;
  reg [31:0] bright_laplace_diff_1_update_0_stage_137;
  reg [31:0] bright_laplace_diff_1_update_0_stage_138;
  reg [31:0] bright_laplace_diff_1_update_0_stage_139;
  reg [31:0] bright_laplace_diff_1_update_0_stage_140;
  reg [31:0] bright_laplace_diff_1_update_0_stage_141;
  reg [31:0] bright_laplace_diff_1_update_0_stage_142;
  reg [31:0] bright_laplace_diff_1_update_0_stage_143;
  reg [31:0] bright_laplace_diff_1_update_0_stage_144;
  reg [31:0] bright_laplace_diff_1_update_0_stage_145;
  reg [31:0] bright_laplace_diff_1_update_0_stage_146;
  reg [31:0] bright_laplace_diff_1_update_0_stage_147;
  reg [31:0] bright_laplace_diff_1_update_0_stage_148;
  reg [31:0] bright_laplace_diff_1_update_0_stage_149;
  reg [31:0] bright_laplace_diff_1_update_0_stage_150;
  reg [31:0] bright_laplace_diff_1_update_0_stage_151;
  reg [31:0] bright_laplace_diff_1_update_0_stage_152;
  reg [31:0] bright_laplace_diff_1_update_0_stage_153;
  reg [31:0] bright_laplace_diff_1_update_0_stage_154;
  reg [31:0] bright_laplace_diff_1_update_0_stage_155;
  reg [31:0] bright_laplace_diff_1_update_0_stage_156;
  reg [31:0] bright_laplace_diff_1_update_0_stage_157;
  reg [31:0] bright_laplace_diff_1_update_0_stage_158;
  reg [31:0] bright_laplace_diff_1_update_0_stage_159;
  reg [31:0] bright_laplace_diff_1_update_0_stage_160;
  reg [31:0] bright_laplace_diff_1_update_0_stage_161;
  reg [31:0] bright_laplace_diff_1_update_0_stage_162;
  reg [31:0] bright_laplace_diff_1_update_0_stage_163;
  reg [31:0] bright_laplace_diff_1_update_0_stage_164;
  reg [31:0] bright_laplace_diff_1_update_0_stage_165;
  reg [31:0] bright_laplace_diff_1_update_0_stage_166;
  reg [31:0] bright_laplace_diff_1_update_0_stage_167;
  reg [31:0] bright_laplace_diff_1_update_0_stage_168;
  reg [31:0] bright_laplace_diff_1_update_0_stage_169;
  reg [31:0] bright_laplace_diff_1_update_0_stage_170;
  reg [31:0] bright_laplace_diff_1_update_0_stage_171;
  reg [31:0] bright_laplace_diff_1_update_0_stage_172;
  reg [31:0] bright_laplace_diff_1_update_0_stage_173;
  reg [31:0] bright_laplace_diff_1_update_0_stage_174;
  reg [31:0] bright_laplace_diff_1_update_0_stage_175;
  reg [31:0] bright_laplace_diff_1_update_0_stage_176;
  reg [31:0] bright_laplace_diff_1_update_0_stage_177;
  reg [31:0] bright_laplace_diff_1_update_0_stage_178;
  reg [31:0] bright_laplace_diff_1_update_0_stage_179;
  reg [31:0] bright_laplace_diff_1_update_0_stage_180;
  reg [31:0] bright_laplace_diff_1_update_0_stage_181;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_103;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_104;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_105;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_106;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_107;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_108;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_109;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_110;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_111;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_112;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_113;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_114;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_115;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_116;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_117;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_118;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_119;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_120;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_121;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_122;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_123;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_124;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_125;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_126;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_127;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_128;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_129;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_130;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_131;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_132;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_133;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_134;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_135;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_136;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_137;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_138;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_139;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_140;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_141;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_142;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_143;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_144;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_145;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_146;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_147;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_148;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_149;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_150;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_151;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_152;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_153;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_154;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_155;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_156;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_157;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_158;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_159;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_160;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_161;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_162;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_163;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_164;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_165;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_166;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_167;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_168;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_169;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_170;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_171;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_172;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_173;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_174;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_175;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_176;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_177;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_178;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_179;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_180;
  reg [31:0] bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_108;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_3_update_0_stage_181;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_109;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_110;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_111;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_112;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_113;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_114;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_115;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_116;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_117;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_118;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_119;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_120;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_121;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_122;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_123;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_124;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_125;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_126;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_127;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_128;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_129;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_130;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_131;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_132;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_133;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_134;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_135;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_136;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_137;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_138;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_139;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_140;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_141;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_142;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_143;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_144;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_145;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_146;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_147;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_148;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_149;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_150;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_151;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_152;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_153;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_154;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_155;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_156;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_157;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_158;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_159;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_160;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_161;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_162;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_163;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_164;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_165;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_166;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_167;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_168;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_169;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_170;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_171;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_172;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_173;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_174;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_175;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_176;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_177;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_178;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_179;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_180;
  reg [31:0] dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_181;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_110;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_111;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_112;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_113;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_114;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_115;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_116;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_117;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_118;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_119;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_120;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_121;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_122;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_123;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_124;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_125;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_126;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_127;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_128;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_129;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_130;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_131;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_132;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_133;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_134;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_135;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_136;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_137;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_138;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_139;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_140;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_141;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_142;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_143;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_144;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_145;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_146;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_147;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_148;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_149;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_150;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_151;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_152;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_153;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_154;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_155;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_156;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_157;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_158;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_159;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_160;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_161;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_162;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_163;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_164;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_165;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_166;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_167;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_168;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_169;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_170;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_171;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_172;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_173;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_174;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_175;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_176;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_177;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_178;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_179;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_180;
  reg [31:0] dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_181;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_111;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_112;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_113;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_114;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_115;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_116;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_117;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_118;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_119;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_120;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_121;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_122;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_123;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_124;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_125;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_126;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_127;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_128;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_129;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_130;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_131;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_132;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_133;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_134;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_135;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_136;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_137;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_138;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_139;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_140;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_141;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_142;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_143;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_144;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_145;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_146;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_147;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_148;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_149;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_150;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_151;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_152;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_153;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_154;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_155;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_156;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_157;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_158;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_159;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_160;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_161;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_162;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_163;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_164;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_165;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_166;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_167;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_168;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_169;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_170;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_171;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_172;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_173;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_174;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_175;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_176;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_177;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_178;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_179;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_180;
  reg [31:0] dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_181;
  reg [31:0] dark_laplace_diff_1_update_0_stage_112;
  reg [31:0] dark_laplace_diff_1_update_0_stage_113;
  reg [31:0] dark_laplace_diff_1_update_0_stage_114;
  reg [31:0] dark_laplace_diff_1_update_0_stage_115;
  reg [31:0] dark_laplace_diff_1_update_0_stage_116;
  reg [31:0] dark_laplace_diff_1_update_0_stage_117;
  reg [31:0] dark_laplace_diff_1_update_0_stage_118;
  reg [31:0] dark_laplace_diff_1_update_0_stage_119;
  reg [31:0] dark_laplace_diff_1_update_0_stage_120;
  reg [31:0] dark_laplace_diff_1_update_0_stage_121;
  reg [31:0] dark_laplace_diff_1_update_0_stage_122;
  reg [31:0] dark_laplace_diff_1_update_0_stage_123;
  reg [31:0] dark_laplace_diff_1_update_0_stage_124;
  reg [31:0] dark_laplace_diff_1_update_0_stage_125;
  reg [31:0] dark_laplace_diff_1_update_0_stage_126;
  reg [31:0] dark_laplace_diff_1_update_0_stage_127;
  reg [31:0] dark_laplace_diff_1_update_0_stage_128;
  reg [31:0] dark_laplace_diff_1_update_0_stage_129;
  reg [31:0] dark_laplace_diff_1_update_0_stage_130;
  reg [31:0] dark_laplace_diff_1_update_0_stage_131;
  reg [31:0] dark_laplace_diff_1_update_0_stage_132;
  reg [31:0] dark_laplace_diff_1_update_0_stage_133;
  reg [31:0] dark_laplace_diff_1_update_0_stage_134;
  reg [31:0] dark_laplace_diff_1_update_0_stage_135;
  reg [31:0] dark_laplace_diff_1_update_0_stage_136;
  reg [31:0] dark_laplace_diff_1_update_0_stage_137;
  reg [31:0] dark_laplace_diff_1_update_0_stage_138;
  reg [31:0] dark_laplace_diff_1_update_0_stage_139;
  reg [31:0] dark_laplace_diff_1_update_0_stage_140;
  reg [31:0] dark_laplace_diff_1_update_0_stage_141;
  reg [31:0] dark_laplace_diff_1_update_0_stage_142;
  reg [31:0] dark_laplace_diff_1_update_0_stage_143;
  reg [31:0] dark_laplace_diff_1_update_0_stage_144;
  reg [31:0] dark_laplace_diff_1_update_0_stage_145;
  reg [31:0] dark_laplace_diff_1_update_0_stage_146;
  reg [31:0] dark_laplace_diff_1_update_0_stage_147;
  reg [31:0] dark_laplace_diff_1_update_0_stage_148;
  reg [31:0] dark_laplace_diff_1_update_0_stage_149;
  reg [31:0] dark_laplace_diff_1_update_0_stage_150;
  reg [31:0] dark_laplace_diff_1_update_0_stage_151;
  reg [31:0] dark_laplace_diff_1_update_0_stage_152;
  reg [31:0] dark_laplace_diff_1_update_0_stage_153;
  reg [31:0] dark_laplace_diff_1_update_0_stage_154;
  reg [31:0] dark_laplace_diff_1_update_0_stage_155;
  reg [31:0] dark_laplace_diff_1_update_0_stage_156;
  reg [31:0] dark_laplace_diff_1_update_0_stage_157;
  reg [31:0] dark_laplace_diff_1_update_0_stage_158;
  reg [31:0] dark_laplace_diff_1_update_0_stage_159;
  reg [31:0] dark_laplace_diff_1_update_0_stage_160;
  reg [31:0] dark_laplace_diff_1_update_0_stage_161;
  reg [31:0] dark_laplace_diff_1_update_0_stage_162;
  reg [31:0] dark_laplace_diff_1_update_0_stage_163;
  reg [31:0] dark_laplace_diff_1_update_0_stage_164;
  reg [31:0] dark_laplace_diff_1_update_0_stage_165;
  reg [31:0] dark_laplace_diff_1_update_0_stage_166;
  reg [31:0] dark_laplace_diff_1_update_0_stage_167;
  reg [31:0] dark_laplace_diff_1_update_0_stage_168;
  reg [31:0] dark_laplace_diff_1_update_0_stage_169;
  reg [31:0] dark_laplace_diff_1_update_0_stage_170;
  reg [31:0] dark_laplace_diff_1_update_0_stage_171;
  reg [31:0] dark_laplace_diff_1_update_0_stage_172;
  reg [31:0] dark_laplace_diff_1_update_0_stage_173;
  reg [31:0] dark_laplace_diff_1_update_0_stage_174;
  reg [31:0] dark_laplace_diff_1_update_0_stage_175;
  reg [31:0] dark_laplace_diff_1_update_0_stage_176;
  reg [31:0] dark_laplace_diff_1_update_0_stage_177;
  reg [31:0] dark_laplace_diff_1_update_0_stage_178;
  reg [31:0] dark_laplace_diff_1_update_0_stage_179;
  reg [31:0] dark_laplace_diff_1_update_0_stage_180;
  reg [31:0] dark_laplace_diff_1_update_0_stage_181;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_113;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_114;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_115;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_116;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_117;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_118;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_119;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_120;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_121;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_122;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_123;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_124;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_125;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_126;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_127;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_128;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_129;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_130;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_131;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_132;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_133;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_134;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_135;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_136;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_137;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_138;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_139;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_140;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_141;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_142;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_143;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_144;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_145;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_146;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_147;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_148;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_149;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_150;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_151;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_152;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_153;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_154;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_155;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_156;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_157;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_158;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_159;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_160;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_161;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_162;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_163;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_164;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_165;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_166;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_167;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_168;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_169;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_170;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_171;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_172;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_173;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_174;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_175;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_176;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_177;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_178;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_179;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_180;
  reg [31:0] dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_181;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_120;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_121;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_122;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_123;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_124;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_125;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_126;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_127;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_128;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_129;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_130;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_131;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_132;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_133;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_134;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_135;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_136;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_137;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_138;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_139;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_140;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_141;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_142;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_143;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_144;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_145;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_146;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_147;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_148;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_149;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_150;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_151;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_152;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_153;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_154;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_155;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_156;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_157;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_158;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_159;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_160;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_161;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_162;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_163;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_164;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_165;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_166;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_167;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_168;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_169;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_170;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_171;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_172;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_173;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_174;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_175;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_176;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_177;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_178;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_179;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_180;
  reg [31:0] bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_181;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_114;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_115;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_116;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_117;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_118;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_119;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_120;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_121;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_122;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_123;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_124;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_125;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_126;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_127;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_128;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_129;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_130;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_131;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_132;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_133;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_134;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_135;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_136;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_137;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_138;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_139;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_140;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_141;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_142;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_143;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_144;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_145;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_146;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_147;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_148;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_149;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_150;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_151;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_152;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_153;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_154;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_155;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_156;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_157;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_158;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_159;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_160;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_161;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_162;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_163;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_164;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_165;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_166;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_167;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_168;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_169;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_170;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_171;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_172;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_173;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_174;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_175;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_176;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_177;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_178;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_179;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_180;
  reg [31:0] bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_181;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_115;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_116;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_117;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_118;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_119;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_120;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_121;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_122;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_123;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_124;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_125;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_126;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_127;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_128;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_129;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_130;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_131;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_132;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_133;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_134;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_135;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_136;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_137;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_138;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_139;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_140;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_141;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_142;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_143;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_144;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_145;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_146;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_147;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_148;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_149;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_150;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_151;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_152;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_153;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_154;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_155;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_156;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_157;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_158;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_159;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_160;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_161;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_162;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_163;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_164;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_165;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_166;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_167;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_168;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_169;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_170;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_171;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_172;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_173;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_174;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_175;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_176;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_177;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_178;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_179;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_180;
  reg [31:0] dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_181;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_116;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_117;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_118;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_119;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_120;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_121;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_122;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_123;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_124;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_125;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_126;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_127;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_128;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_129;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_130;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_131;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_132;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_133;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_134;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_135;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_136;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_137;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_138;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_139;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_140;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_141;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_142;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_143;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_144;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_145;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_146;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_147;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_148;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_149;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_150;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_151;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_152;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_153;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_154;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_155;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_156;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_157;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_158;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_159;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_160;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_161;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_162;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_163;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_164;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_165;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_166;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_167;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_168;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_169;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_170;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_171;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_172;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_173;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_174;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_175;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_176;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_177;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_178;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_179;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_180;
  reg [31:0] bright_weights_normed_fused_level_0_update_0_read_read_79_stage_181;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_117;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_118;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_119;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_120;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_121;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_122;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_123;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_124;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_125;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_126;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_127;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_128;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_129;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_130;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_131;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_132;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_133;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_134;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_135;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_136;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_137;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_138;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_139;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_140;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_141;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_142;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_143;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_144;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_145;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_146;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_147;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_148;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_149;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_150;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_151;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_152;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_153;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_154;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_155;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_156;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_157;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_158;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_159;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_160;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_161;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_162;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_163;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_164;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_165;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_166;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_167;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_168;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_169;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_170;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_171;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_172;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_173;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_174;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_175;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_176;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_177;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_178;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_179;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_180;
  reg [31:0] dark_weights_normed_fused_level_0_update_0_read_read_80_stage_181;
  reg [31:0] fused_level_0_update_0_stage_118;
  reg [31:0] fused_level_0_update_0_stage_119;
  reg [31:0] fused_level_0_update_0_stage_120;
  reg [31:0] fused_level_0_update_0_stage_121;
  reg [31:0] fused_level_0_update_0_stage_122;
  reg [31:0] fused_level_0_update_0_stage_123;
  reg [31:0] fused_level_0_update_0_stage_124;
  reg [31:0] fused_level_0_update_0_stage_125;
  reg [31:0] fused_level_0_update_0_stage_126;
  reg [31:0] fused_level_0_update_0_stage_127;
  reg [31:0] fused_level_0_update_0_stage_128;
  reg [31:0] fused_level_0_update_0_stage_129;
  reg [31:0] fused_level_0_update_0_stage_130;
  reg [31:0] fused_level_0_update_0_stage_131;
  reg [31:0] fused_level_0_update_0_stage_132;
  reg [31:0] fused_level_0_update_0_stage_133;
  reg [31:0] fused_level_0_update_0_stage_134;
  reg [31:0] fused_level_0_update_0_stage_135;
  reg [31:0] fused_level_0_update_0_stage_136;
  reg [31:0] fused_level_0_update_0_stage_137;
  reg [31:0] fused_level_0_update_0_stage_138;
  reg [31:0] fused_level_0_update_0_stage_139;
  reg [31:0] fused_level_0_update_0_stage_140;
  reg [31:0] fused_level_0_update_0_stage_141;
  reg [31:0] fused_level_0_update_0_stage_142;
  reg [31:0] fused_level_0_update_0_stage_143;
  reg [31:0] fused_level_0_update_0_stage_144;
  reg [31:0] fused_level_0_update_0_stage_145;
  reg [31:0] fused_level_0_update_0_stage_146;
  reg [31:0] fused_level_0_update_0_stage_147;
  reg [31:0] fused_level_0_update_0_stage_148;
  reg [31:0] fused_level_0_update_0_stage_149;
  reg [31:0] fused_level_0_update_0_stage_150;
  reg [31:0] fused_level_0_update_0_stage_151;
  reg [31:0] fused_level_0_update_0_stage_152;
  reg [31:0] fused_level_0_update_0_stage_153;
  reg [31:0] fused_level_0_update_0_stage_154;
  reg [31:0] fused_level_0_update_0_stage_155;
  reg [31:0] fused_level_0_update_0_stage_156;
  reg [31:0] fused_level_0_update_0_stage_157;
  reg [31:0] fused_level_0_update_0_stage_158;
  reg [31:0] fused_level_0_update_0_stage_159;
  reg [31:0] fused_level_0_update_0_stage_160;
  reg [31:0] fused_level_0_update_0_stage_161;
  reg [31:0] fused_level_0_update_0_stage_162;
  reg [31:0] fused_level_0_update_0_stage_163;
  reg [31:0] fused_level_0_update_0_stage_164;
  reg [31:0] fused_level_0_update_0_stage_165;
  reg [31:0] fused_level_0_update_0_stage_166;
  reg [31:0] fused_level_0_update_0_stage_167;
  reg [31:0] fused_level_0_update_0_stage_168;
  reg [31:0] fused_level_0_update_0_stage_169;
  reg [31:0] fused_level_0_update_0_stage_170;
  reg [31:0] fused_level_0_update_0_stage_171;
  reg [31:0] fused_level_0_update_0_stage_172;
  reg [31:0] fused_level_0_update_0_stage_173;
  reg [31:0] fused_level_0_update_0_stage_174;
  reg [31:0] fused_level_0_update_0_stage_175;
  reg [31:0] fused_level_0_update_0_stage_176;
  reg [31:0] fused_level_0_update_0_stage_177;
  reg [31:0] fused_level_0_update_0_stage_178;
  reg [31:0] fused_level_0_update_0_stage_179;
  reg [31:0] fused_level_0_update_0_stage_180;
  reg [31:0] fused_level_0_update_0_stage_181;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_119;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_120;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_121;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_122;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_123;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_124;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_125;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_126;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_127;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_128;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_129;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_130;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_131;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_132;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_133;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_134;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_135;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_136;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_137;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_138;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_139;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_140;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_141;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_142;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_143;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_144;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_145;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_146;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_147;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_148;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_149;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_150;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_151;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_152;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_153;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_154;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_155;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_156;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_157;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_158;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_159;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_160;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_161;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_162;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_163;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_164;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_165;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_166;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_167;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_168;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_169;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_170;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_171;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_172;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_173;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_174;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_175;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_176;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_177;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_178;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_179;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_180;
  reg [31:0] fused_level_0_fused_level_0_update_0_write_write_81_stage_181;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_121;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_122;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_123;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_124;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_125;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_126;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_127;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_128;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_129;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_130;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_131;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_132;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_133;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_134;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_135;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_136;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_137;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_138;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_139;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_140;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_141;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_142;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_143;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_144;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_145;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_146;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_147;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_148;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_149;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_150;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_151;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_152;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_153;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_154;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_155;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_156;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_157;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_158;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_159;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_160;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_161;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_162;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_163;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_164;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_165;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_166;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_167;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_168;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_169;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_170;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_171;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_172;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_173;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_174;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_175;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_176;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_177;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_178;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_179;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_180;
  reg [31:0] bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_181;
  reg [31:0] bright_laplace_diff_2_update_0_stage_122;
  reg [31:0] bright_laplace_diff_2_update_0_stage_123;
  reg [31:0] bright_laplace_diff_2_update_0_stage_124;
  reg [31:0] bright_laplace_diff_2_update_0_stage_125;
  reg [31:0] bright_laplace_diff_2_update_0_stage_126;
  reg [31:0] bright_laplace_diff_2_update_0_stage_127;
  reg [31:0] bright_laplace_diff_2_update_0_stage_128;
  reg [31:0] bright_laplace_diff_2_update_0_stage_129;
  reg [31:0] bright_laplace_diff_2_update_0_stage_130;
  reg [31:0] bright_laplace_diff_2_update_0_stage_131;
  reg [31:0] bright_laplace_diff_2_update_0_stage_132;
  reg [31:0] bright_laplace_diff_2_update_0_stage_133;
  reg [31:0] bright_laplace_diff_2_update_0_stage_134;
  reg [31:0] bright_laplace_diff_2_update_0_stage_135;
  reg [31:0] bright_laplace_diff_2_update_0_stage_136;
  reg [31:0] bright_laplace_diff_2_update_0_stage_137;
  reg [31:0] bright_laplace_diff_2_update_0_stage_138;
  reg [31:0] bright_laplace_diff_2_update_0_stage_139;
  reg [31:0] bright_laplace_diff_2_update_0_stage_140;
  reg [31:0] bright_laplace_diff_2_update_0_stage_141;
  reg [31:0] bright_laplace_diff_2_update_0_stage_142;
  reg [31:0] bright_laplace_diff_2_update_0_stage_143;
  reg [31:0] bright_laplace_diff_2_update_0_stage_144;
  reg [31:0] bright_laplace_diff_2_update_0_stage_145;
  reg [31:0] bright_laplace_diff_2_update_0_stage_146;
  reg [31:0] bright_laplace_diff_2_update_0_stage_147;
  reg [31:0] bright_laplace_diff_2_update_0_stage_148;
  reg [31:0] bright_laplace_diff_2_update_0_stage_149;
  reg [31:0] bright_laplace_diff_2_update_0_stage_150;
  reg [31:0] bright_laplace_diff_2_update_0_stage_151;
  reg [31:0] bright_laplace_diff_2_update_0_stage_152;
  reg [31:0] bright_laplace_diff_2_update_0_stage_153;
  reg [31:0] bright_laplace_diff_2_update_0_stage_154;
  reg [31:0] bright_laplace_diff_2_update_0_stage_155;
  reg [31:0] bright_laplace_diff_2_update_0_stage_156;
  reg [31:0] bright_laplace_diff_2_update_0_stage_157;
  reg [31:0] bright_laplace_diff_2_update_0_stage_158;
  reg [31:0] bright_laplace_diff_2_update_0_stage_159;
  reg [31:0] bright_laplace_diff_2_update_0_stage_160;
  reg [31:0] bright_laplace_diff_2_update_0_stage_161;
  reg [31:0] bright_laplace_diff_2_update_0_stage_162;
  reg [31:0] bright_laplace_diff_2_update_0_stage_163;
  reg [31:0] bright_laplace_diff_2_update_0_stage_164;
  reg [31:0] bright_laplace_diff_2_update_0_stage_165;
  reg [31:0] bright_laplace_diff_2_update_0_stage_166;
  reg [31:0] bright_laplace_diff_2_update_0_stage_167;
  reg [31:0] bright_laplace_diff_2_update_0_stage_168;
  reg [31:0] bright_laplace_diff_2_update_0_stage_169;
  reg [31:0] bright_laplace_diff_2_update_0_stage_170;
  reg [31:0] bright_laplace_diff_2_update_0_stage_171;
  reg [31:0] bright_laplace_diff_2_update_0_stage_172;
  reg [31:0] bright_laplace_diff_2_update_0_stage_173;
  reg [31:0] bright_laplace_diff_2_update_0_stage_174;
  reg [31:0] bright_laplace_diff_2_update_0_stage_175;
  reg [31:0] bright_laplace_diff_2_update_0_stage_176;
  reg [31:0] bright_laplace_diff_2_update_0_stage_177;
  reg [31:0] bright_laplace_diff_2_update_0_stage_178;
  reg [31:0] bright_laplace_diff_2_update_0_stage_179;
  reg [31:0] bright_laplace_diff_2_update_0_stage_180;
  reg [31:0] bright_laplace_diff_2_update_0_stage_181;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_123;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_124;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_125;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_126;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_127;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_128;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_129;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_130;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_131;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_132;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_133;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_134;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_135;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_136;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_137;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_138;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_139;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_140;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_141;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_142;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_143;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_144;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_145;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_146;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_147;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_148;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_149;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_150;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_151;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_152;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_153;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_154;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_155;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_156;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_157;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_158;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_159;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_160;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_161;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_162;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_163;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_164;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_165;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_166;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_167;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_168;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_169;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_170;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_171;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_172;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_173;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_174;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_175;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_176;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_177;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_178;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_179;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_180;
  reg [31:0] bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_181;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_130;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_131;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_132;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_133;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_134;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_135;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_136;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_137;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_138;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_139;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_140;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_141;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_142;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_143;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_144;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_145;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_146;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_147;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_148;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_149;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_150;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_151;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_152;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_153;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_154;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_155;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_156;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_157;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_158;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_159;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_160;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_161;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_162;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_163;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_164;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_165;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_166;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_167;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_168;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_169;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_170;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_171;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_172;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_173;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_174;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_175;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_176;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_177;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_178;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_179;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_180;
  reg [287:0] bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_181;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_124;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_125;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_126;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_127;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_128;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_129;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_130;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_131;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_132;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_133;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_134;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_135;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_136;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_137;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_138;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_139;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_140;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_141;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_142;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_143;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_144;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_145;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_146;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_147;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_148;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_149;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_150;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_151;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_152;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_153;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_154;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_155;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_156;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_157;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_158;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_159;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_160;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_161;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_162;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_163;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_164;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_165;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_166;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_167;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_168;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_169;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_170;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_171;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_172;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_173;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_174;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_175;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_176;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_177;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_178;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_179;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_180;
  reg [31:0] bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_181;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_125;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_126;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_127;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_128;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_129;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_130;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_131;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_132;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_133;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_134;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_135;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_136;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_137;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_138;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_139;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_140;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_141;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_142;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_143;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_144;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_145;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_146;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_147;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_148;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_149;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_150;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_151;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_152;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_153;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_154;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_155;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_156;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_157;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_158;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_159;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_160;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_161;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_162;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_163;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_164;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_165;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_166;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_167;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_168;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_169;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_170;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_171;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_172;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_173;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_174;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_175;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_176;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_177;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_178;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_179;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_180;
  reg [31:0] dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_131;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_132;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_133;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_134;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_135;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_136;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_137;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_138;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_2_update_0_stage_181;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_133;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_134;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_135;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_136;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_137;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_138;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_139;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_140;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_141;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_142;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_143;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_144;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_145;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_146;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_147;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_148;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_149;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_150;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_151;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_152;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_153;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_154;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_155;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_156;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_157;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_158;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_159;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_160;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_161;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_162;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_163;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_164;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_165;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_166;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_167;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_168;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_169;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_170;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_171;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_172;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_173;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_174;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_175;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_176;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_177;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_178;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_179;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_180;
  reg [31:0] dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_132;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_133;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_134;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_135;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_136;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_137;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_138;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_181;
  reg [31:0] dark_gauss_ds_3_update_0_stage_134;
  reg [31:0] dark_gauss_ds_3_update_0_stage_135;
  reg [31:0] dark_gauss_ds_3_update_0_stage_136;
  reg [31:0] dark_gauss_ds_3_update_0_stage_137;
  reg [31:0] dark_gauss_ds_3_update_0_stage_138;
  reg [31:0] dark_gauss_ds_3_update_0_stage_139;
  reg [31:0] dark_gauss_ds_3_update_0_stage_140;
  reg [31:0] dark_gauss_ds_3_update_0_stage_141;
  reg [31:0] dark_gauss_ds_3_update_0_stage_142;
  reg [31:0] dark_gauss_ds_3_update_0_stage_143;
  reg [31:0] dark_gauss_ds_3_update_0_stage_144;
  reg [31:0] dark_gauss_ds_3_update_0_stage_145;
  reg [31:0] dark_gauss_ds_3_update_0_stage_146;
  reg [31:0] dark_gauss_ds_3_update_0_stage_147;
  reg [31:0] dark_gauss_ds_3_update_0_stage_148;
  reg [31:0] dark_gauss_ds_3_update_0_stage_149;
  reg [31:0] dark_gauss_ds_3_update_0_stage_150;
  reg [31:0] dark_gauss_ds_3_update_0_stage_151;
  reg [31:0] dark_gauss_ds_3_update_0_stage_152;
  reg [31:0] dark_gauss_ds_3_update_0_stage_153;
  reg [31:0] dark_gauss_ds_3_update_0_stage_154;
  reg [31:0] dark_gauss_ds_3_update_0_stage_155;
  reg [31:0] dark_gauss_ds_3_update_0_stage_156;
  reg [31:0] dark_gauss_ds_3_update_0_stage_157;
  reg [31:0] dark_gauss_ds_3_update_0_stage_158;
  reg [31:0] dark_gauss_ds_3_update_0_stage_159;
  reg [31:0] dark_gauss_ds_3_update_0_stage_160;
  reg [31:0] dark_gauss_ds_3_update_0_stage_161;
  reg [31:0] dark_gauss_ds_3_update_0_stage_162;
  reg [31:0] dark_gauss_ds_3_update_0_stage_163;
  reg [31:0] dark_gauss_ds_3_update_0_stage_164;
  reg [31:0] dark_gauss_ds_3_update_0_stage_165;
  reg [31:0] dark_gauss_ds_3_update_0_stage_166;
  reg [31:0] dark_gauss_ds_3_update_0_stage_167;
  reg [31:0] dark_gauss_ds_3_update_0_stage_168;
  reg [31:0] dark_gauss_ds_3_update_0_stage_169;
  reg [31:0] dark_gauss_ds_3_update_0_stage_170;
  reg [31:0] dark_gauss_ds_3_update_0_stage_171;
  reg [31:0] dark_gauss_ds_3_update_0_stage_172;
  reg [31:0] dark_gauss_ds_3_update_0_stage_173;
  reg [31:0] dark_gauss_ds_3_update_0_stage_174;
  reg [31:0] dark_gauss_ds_3_update_0_stage_175;
  reg [31:0] dark_gauss_ds_3_update_0_stage_176;
  reg [31:0] dark_gauss_ds_3_update_0_stage_177;
  reg [31:0] dark_gauss_ds_3_update_0_stage_178;
  reg [31:0] dark_gauss_ds_3_update_0_stage_179;
  reg [31:0] dark_gauss_ds_3_update_0_stage_180;
  reg [31:0] dark_gauss_ds_3_update_0_stage_181;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_135;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_136;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_137;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_138;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_139;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_140;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_141;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_142;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_143;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_144;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_145;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_146;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_147;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_148;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_149;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_150;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_151;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_152;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_153;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_154;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_155;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_156;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_157;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_158;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_159;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_160;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_161;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_162;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_163;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_164;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_165;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_166;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_167;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_168;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_169;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_170;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_171;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_172;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_173;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_174;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_175;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_176;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_177;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_178;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_179;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_180;
  reg [31:0] dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_139;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_140;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_141;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_142;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_143;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_144;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_145;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_146;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_147;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_148;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_149;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_140;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_141;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_142;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_143;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_144;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_145;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_146;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_147;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_148;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_149;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_150;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_151;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_152;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_2_update_0_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_141;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_142;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_143;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_144;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_145;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_146;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_147;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_148;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_149;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_150;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_151;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_152;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_181;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_145;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_146;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_147;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_148;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_149;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_150;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_151;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_152;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_153;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_154;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_155;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_156;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_157;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_158;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_159;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_160;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_161;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_162;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_163;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_164;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_165;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_166;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_167;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_168;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_169;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_170;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_171;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_172;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_173;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_174;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_175;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_176;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_177;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_178;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_179;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_180;
  reg [31:0] dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_181;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_146;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_147;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_148;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_149;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_150;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_151;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_152;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_153;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_154;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_155;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_156;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_157;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_158;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_159;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_160;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_161;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_162;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_163;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_164;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_165;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_166;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_167;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_168;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_169;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_170;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_171;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_172;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_173;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_174;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_175;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_176;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_177;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_178;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_179;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_180;
  reg [31:0] dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_181;
  reg [31:0] dark_laplace_diff_2_update_0_stage_147;
  reg [31:0] dark_laplace_diff_2_update_0_stage_148;
  reg [31:0] dark_laplace_diff_2_update_0_stage_149;
  reg [31:0] dark_laplace_diff_2_update_0_stage_150;
  reg [31:0] dark_laplace_diff_2_update_0_stage_151;
  reg [31:0] dark_laplace_diff_2_update_0_stage_152;
  reg [31:0] dark_laplace_diff_2_update_0_stage_153;
  reg [31:0] dark_laplace_diff_2_update_0_stage_154;
  reg [31:0] dark_laplace_diff_2_update_0_stage_155;
  reg [31:0] dark_laplace_diff_2_update_0_stage_156;
  reg [31:0] dark_laplace_diff_2_update_0_stage_157;
  reg [31:0] dark_laplace_diff_2_update_0_stage_158;
  reg [31:0] dark_laplace_diff_2_update_0_stage_159;
  reg [31:0] dark_laplace_diff_2_update_0_stage_160;
  reg [31:0] dark_laplace_diff_2_update_0_stage_161;
  reg [31:0] dark_laplace_diff_2_update_0_stage_162;
  reg [31:0] dark_laplace_diff_2_update_0_stage_163;
  reg [31:0] dark_laplace_diff_2_update_0_stage_164;
  reg [31:0] dark_laplace_diff_2_update_0_stage_165;
  reg [31:0] dark_laplace_diff_2_update_0_stage_166;
  reg [31:0] dark_laplace_diff_2_update_0_stage_167;
  reg [31:0] dark_laplace_diff_2_update_0_stage_168;
  reg [31:0] dark_laplace_diff_2_update_0_stage_169;
  reg [31:0] dark_laplace_diff_2_update_0_stage_170;
  reg [31:0] dark_laplace_diff_2_update_0_stage_171;
  reg [31:0] dark_laplace_diff_2_update_0_stage_172;
  reg [31:0] dark_laplace_diff_2_update_0_stage_173;
  reg [31:0] dark_laplace_diff_2_update_0_stage_174;
  reg [31:0] dark_laplace_diff_2_update_0_stage_175;
  reg [31:0] dark_laplace_diff_2_update_0_stage_176;
  reg [31:0] dark_laplace_diff_2_update_0_stage_177;
  reg [31:0] dark_laplace_diff_2_update_0_stage_178;
  reg [31:0] dark_laplace_diff_2_update_0_stage_179;
  reg [31:0] dark_laplace_diff_2_update_0_stage_180;
  reg [31:0] dark_laplace_diff_2_update_0_stage_181;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_149;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_150;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_151;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_152;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_153;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_154;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_155;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_156;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_157;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_158;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_159;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_160;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_161;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_162;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_163;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_164;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_165;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_166;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_167;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_168;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_169;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_170;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_171;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_172;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_173;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_174;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_175;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_176;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_177;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_178;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_179;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_180;
  reg [287:0] bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_150;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_3_update_0_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_151;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_181;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_152;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_153;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_154;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_155;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_156;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_157;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_158;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_159;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_160;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_161;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_162;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_163;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_164;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_165;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_166;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_167;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_168;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_169;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_170;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_171;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_172;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_173;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_174;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_175;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_176;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_177;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_178;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_179;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_180;
  reg [31:0] bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_153;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_3_update_0_stage_181;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_155;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_156;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_157;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_158;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_159;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_160;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_161;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_162;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_163;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_164;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_165;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_166;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_167;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_168;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_169;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_170;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_171;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_172;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_173;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_174;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_175;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_176;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_177;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_178;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_179;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_180;
  reg [31:0] bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_154;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_155;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_156;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_181;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_156;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_157;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_158;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_159;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_160;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_161;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_162;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_163;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_164;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_165;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_166;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_167;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_168;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_169;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_170;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_171;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_172;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_173;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_174;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_175;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_176;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_177;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_178;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_179;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_180;
  reg [31:0] dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_181;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_157;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_158;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_159;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_160;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_161;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_162;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_163;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_164;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_165;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_166;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_167;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_168;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_169;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_170;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_171;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_172;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_173;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_174;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_175;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_176;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_177;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_178;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_179;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_180;
  reg [31:0] bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_181;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_158;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_159;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_160;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_161;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_162;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_163;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_164;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_165;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_166;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_167;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_168;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_169;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_170;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_171;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_172;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_173;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_174;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_175;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_176;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_177;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_178;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_179;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_180;
  reg [31:0] dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_181;
  reg [31:0] fused_level_2_update_0_stage_159;
  reg [31:0] fused_level_2_update_0_stage_160;
  reg [31:0] fused_level_2_update_0_stage_161;
  reg [31:0] fused_level_2_update_0_stage_162;
  reg [31:0] fused_level_2_update_0_stage_163;
  reg [31:0] fused_level_2_update_0_stage_164;
  reg [31:0] fused_level_2_update_0_stage_165;
  reg [31:0] fused_level_2_update_0_stage_166;
  reg [31:0] fused_level_2_update_0_stage_167;
  reg [31:0] fused_level_2_update_0_stage_168;
  reg [31:0] fused_level_2_update_0_stage_169;
  reg [31:0] fused_level_2_update_0_stage_170;
  reg [31:0] fused_level_2_update_0_stage_171;
  reg [31:0] fused_level_2_update_0_stage_172;
  reg [31:0] fused_level_2_update_0_stage_173;
  reg [31:0] fused_level_2_update_0_stage_174;
  reg [31:0] fused_level_2_update_0_stage_175;
  reg [31:0] fused_level_2_update_0_stage_176;
  reg [31:0] fused_level_2_update_0_stage_177;
  reg [31:0] fused_level_2_update_0_stage_178;
  reg [31:0] fused_level_2_update_0_stage_179;
  reg [31:0] fused_level_2_update_0_stage_180;
  reg [31:0] fused_level_2_update_0_stage_181;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_160;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_161;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_162;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_163;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_164;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_165;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_166;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_167;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_168;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_169;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_170;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_171;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_172;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_173;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_174;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_175;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_176;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_177;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_178;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_179;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_180;
  reg [31:0] fused_level_2_fused_level_2_update_0_write_write_111_stage_181;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_161;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_162;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_163;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_164;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_165;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_166;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_167;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_168;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_169;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_170;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_171;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_172;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_173;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_174;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_175;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_176;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_177;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_178;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_179;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_180;
  reg [31:0] bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_181;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_162;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_163;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_164;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_165;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_166;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_167;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_168;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_169;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_170;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_171;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_172;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_173;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_174;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_175;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_176;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_177;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_178;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_179;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_180;
  reg [31:0] dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_181;


  always @(posedge clk) begin
    if (rst) begin
      started <= 0;
      stage_1_active <= 0;
      stage_2_active <= 0;
      stage_3_active <= 0;
      stage_4_active <= 0;
      stage_5_active <= 0;
      stage_6_active <= 0;
      stage_7_active <= 0;
      stage_8_active <= 0;
      stage_9_active <= 0;
      stage_10_active <= 0;
      stage_11_active <= 0;
      stage_12_active <= 0;
      stage_13_active <= 0;
      stage_14_active <= 0;
      stage_15_active <= 0;
      stage_16_active <= 0;
      stage_17_active <= 0;
      stage_18_active <= 0;
      stage_19_active <= 0;
      stage_20_active <= 0;
      stage_21_active <= 0;
      stage_22_active <= 0;
      stage_23_active <= 0;
      stage_24_active <= 0;
      stage_25_active <= 0;
      stage_26_active <= 0;
      stage_27_active <= 0;
      stage_28_active <= 0;
      stage_29_active <= 0;
      stage_30_active <= 0;
      stage_31_active <= 0;
      stage_32_active <= 0;
      stage_33_active <= 0;
      stage_34_active <= 0;
      stage_35_active <= 0;
      stage_36_active <= 0;
      stage_37_active <= 0;
      stage_38_active <= 0;
      stage_39_active <= 0;
      stage_40_active <= 0;
      stage_41_active <= 0;
      stage_42_active <= 0;
      stage_43_active <= 0;
      stage_44_active <= 0;
      stage_45_active <= 0;
      stage_46_active <= 0;
      stage_47_active <= 0;
      stage_48_active <= 0;
      stage_49_active <= 0;
      stage_50_active <= 0;
      stage_51_active <= 0;
      stage_52_active <= 0;
      stage_53_active <= 0;
      stage_54_active <= 0;
      stage_55_active <= 0;
      stage_56_active <= 0;
      stage_57_active <= 0;
      stage_58_active <= 0;
      stage_59_active <= 0;
      stage_60_active <= 0;
      stage_61_active <= 0;
      stage_62_active <= 0;
      stage_63_active <= 0;
      stage_64_active <= 0;
      stage_65_active <= 0;
      stage_66_active <= 0;
      stage_67_active <= 0;
      stage_68_active <= 0;
      stage_69_active <= 0;
      stage_70_active <= 0;
      stage_71_active <= 0;
      stage_72_active <= 0;
      stage_73_active <= 0;
      stage_74_active <= 0;
      stage_75_active <= 0;
      stage_76_active <= 0;
      stage_77_active <= 0;
      stage_78_active <= 0;
      stage_79_active <= 0;
      stage_80_active <= 0;
      stage_81_active <= 0;
      stage_82_active <= 0;
      stage_83_active <= 0;
      stage_84_active <= 0;
      stage_85_active <= 0;
      stage_86_active <= 0;
      stage_87_active <= 0;
      stage_88_active <= 0;
      stage_89_active <= 0;
      stage_90_active <= 0;
      stage_91_active <= 0;
      stage_92_active <= 0;
      stage_93_active <= 0;
      stage_94_active <= 0;
      stage_95_active <= 0;
      stage_96_active <= 0;
      stage_97_active <= 0;
      stage_98_active <= 0;
      stage_99_active <= 0;
      stage_100_active <= 0;
      stage_101_active <= 0;
      stage_102_active <= 0;
      stage_103_active <= 0;
      stage_104_active <= 0;
      stage_105_active <= 0;
      stage_106_active <= 0;
      stage_107_active <= 0;
      stage_108_active <= 0;
      stage_109_active <= 0;
      stage_110_active <= 0;
      stage_111_active <= 0;
      stage_112_active <= 0;
      stage_113_active <= 0;
      stage_114_active <= 0;
      stage_115_active <= 0;
      stage_116_active <= 0;
      stage_117_active <= 0;
      stage_118_active <= 0;
      stage_119_active <= 0;
      stage_120_active <= 0;
      stage_121_active <= 0;
      stage_122_active <= 0;
      stage_123_active <= 0;
      stage_124_active <= 0;
      stage_125_active <= 0;
      stage_126_active <= 0;
      stage_127_active <= 0;
      stage_128_active <= 0;
      stage_129_active <= 0;
      stage_130_active <= 0;
      stage_131_active <= 0;
      stage_132_active <= 0;
      stage_133_active <= 0;
      stage_134_active <= 0;
      stage_135_active <= 0;
      stage_136_active <= 0;
      stage_137_active <= 0;
      stage_138_active <= 0;
      stage_139_active <= 0;
      stage_140_active <= 0;
      stage_141_active <= 0;
      stage_142_active <= 0;
      stage_143_active <= 0;
      stage_144_active <= 0;
      stage_145_active <= 0;
      stage_146_active <= 0;
      stage_147_active <= 0;
      stage_148_active <= 0;
      stage_149_active <= 0;
      stage_150_active <= 0;
      stage_151_active <= 0;
      stage_152_active <= 0;
      stage_153_active <= 0;
      stage_154_active <= 0;
      stage_155_active <= 0;
      stage_156_active <= 0;
      stage_157_active <= 0;
      stage_158_active <= 0;
      stage_159_active <= 0;
      stage_160_active <= 0;
      stage_161_active <= 0;
      stage_162_active <= 0;
      stage_163_active <= 0;
      stage_164_active <= 0;
      stage_165_active <= 0;
      stage_166_active <= 0;
      stage_167_active <= 0;
      stage_168_active <= 0;
      stage_169_active <= 0;
      stage_170_active <= 0;
      stage_171_active <= 0;
      stage_172_active <= 0;
      stage_173_active <= 0;
      stage_174_active <= 0;
      stage_175_active <= 0;
      stage_176_active <= 0;
      stage_177_active <= 0;
      stage_178_active <= 0;
      stage_179_active <= 0;
      stage_180_active <= 0;
    end else begin

      if (start) begin
        started <= 1;
      end

      stage_1_active <= stage_0_active;
      stage_1_at_iter_0 <= stage_0_at_iter_0;
      stage_2_active <= stage_1_active;
      stage_2_at_iter_0 <= stage_1_at_iter_0;
      stage_3_active <= stage_2_active;
      stage_3_at_iter_0 <= stage_2_at_iter_0;
      stage_4_active <= stage_3_active;
      stage_4_at_iter_0 <= stage_3_at_iter_0;
      stage_5_active <= stage_4_active;
      stage_5_at_iter_0 <= stage_4_at_iter_0;
      stage_6_active <= stage_5_active;
      stage_6_at_iter_0 <= stage_5_at_iter_0;
      stage_7_active <= stage_6_active;
      stage_7_at_iter_0 <= stage_6_at_iter_0;
      stage_8_active <= stage_7_active;
      stage_8_at_iter_0 <= stage_7_at_iter_0;
      stage_9_active <= stage_8_active;
      stage_9_at_iter_0 <= stage_8_at_iter_0;
      stage_10_active <= stage_9_active;
      stage_10_at_iter_0 <= stage_9_at_iter_0;
      stage_11_active <= stage_10_active;
      stage_11_at_iter_0 <= stage_10_at_iter_0;
      stage_12_active <= stage_11_active;
      stage_12_at_iter_0 <= stage_11_at_iter_0;
      stage_13_active <= stage_12_active;
      stage_13_at_iter_0 <= stage_12_at_iter_0;
      stage_14_active <= stage_13_active;
      stage_14_at_iter_0 <= stage_13_at_iter_0;
      stage_15_active <= stage_14_active;
      stage_15_at_iter_0 <= stage_14_at_iter_0;
      stage_16_active <= stage_15_active;
      stage_16_at_iter_0 <= stage_15_at_iter_0;
      stage_17_active <= stage_16_active;
      stage_17_at_iter_0 <= stage_16_at_iter_0;
      stage_18_active <= stage_17_active;
      stage_18_at_iter_0 <= stage_17_at_iter_0;
      stage_19_active <= stage_18_active;
      stage_19_at_iter_0 <= stage_18_at_iter_0;
      stage_20_active <= stage_19_active;
      stage_20_at_iter_0 <= stage_19_at_iter_0;
      stage_21_active <= stage_20_active;
      stage_21_at_iter_0 <= stage_20_at_iter_0;
      stage_22_active <= stage_21_active;
      stage_22_at_iter_0 <= stage_21_at_iter_0;
      stage_23_active <= stage_22_active;
      stage_23_at_iter_0 <= stage_22_at_iter_0;
      stage_24_active <= stage_23_active;
      stage_24_at_iter_0 <= stage_23_at_iter_0;
      stage_25_active <= stage_24_active;
      stage_25_at_iter_0 <= stage_24_at_iter_0;
      stage_26_active <= stage_25_active;
      stage_26_at_iter_0 <= stage_25_at_iter_0;
      stage_27_active <= stage_26_active;
      stage_27_at_iter_0 <= stage_26_at_iter_0;
      stage_28_active <= stage_27_active;
      stage_28_at_iter_0 <= stage_27_at_iter_0;
      stage_29_active <= stage_28_active;
      stage_29_at_iter_0 <= stage_28_at_iter_0;
      stage_30_active <= stage_29_active;
      stage_30_at_iter_0 <= stage_29_at_iter_0;
      stage_31_active <= stage_30_active;
      stage_31_at_iter_0 <= stage_30_at_iter_0;
      stage_32_active <= stage_31_active;
      stage_32_at_iter_0 <= stage_31_at_iter_0;
      stage_33_active <= stage_32_active;
      stage_33_at_iter_0 <= stage_32_at_iter_0;
      stage_34_active <= stage_33_active;
      stage_34_at_iter_0 <= stage_33_at_iter_0;
      stage_35_active <= stage_34_active;
      stage_35_at_iter_0 <= stage_34_at_iter_0;
      stage_36_active <= stage_35_active;
      stage_36_at_iter_0 <= stage_35_at_iter_0;
      stage_37_active <= stage_36_active;
      stage_37_at_iter_0 <= stage_36_at_iter_0;
      stage_38_active <= stage_37_active;
      stage_38_at_iter_0 <= stage_37_at_iter_0;
      stage_39_active <= stage_38_active;
      stage_39_at_iter_0 <= stage_38_at_iter_0;
      stage_40_active <= stage_39_active;
      stage_40_at_iter_0 <= stage_39_at_iter_0;
      stage_41_active <= stage_40_active;
      stage_41_at_iter_0 <= stage_40_at_iter_0;
      stage_42_active <= stage_41_active;
      stage_42_at_iter_0 <= stage_41_at_iter_0;
      stage_43_active <= stage_42_active;
      stage_43_at_iter_0 <= stage_42_at_iter_0;
      stage_44_active <= stage_43_active;
      stage_44_at_iter_0 <= stage_43_at_iter_0;
      stage_45_active <= stage_44_active;
      stage_45_at_iter_0 <= stage_44_at_iter_0;
      stage_46_active <= stage_45_active;
      stage_46_at_iter_0 <= stage_45_at_iter_0;
      stage_47_active <= stage_46_active;
      stage_47_at_iter_0 <= stage_46_at_iter_0;
      stage_48_active <= stage_47_active;
      stage_48_at_iter_0 <= stage_47_at_iter_0;
      stage_49_active <= stage_48_active;
      stage_49_at_iter_0 <= stage_48_at_iter_0;
      stage_50_active <= stage_49_active;
      stage_50_at_iter_0 <= stage_49_at_iter_0;
      stage_51_active <= stage_50_active;
      stage_51_at_iter_0 <= stage_50_at_iter_0;
      stage_52_active <= stage_51_active;
      stage_52_at_iter_0 <= stage_51_at_iter_0;
      stage_53_active <= stage_52_active;
      stage_53_at_iter_0 <= stage_52_at_iter_0;
      stage_54_active <= stage_53_active;
      stage_54_at_iter_0 <= stage_53_at_iter_0;
      stage_55_active <= stage_54_active;
      stage_55_at_iter_0 <= stage_54_at_iter_0;
      stage_56_active <= stage_55_active;
      stage_56_at_iter_0 <= stage_55_at_iter_0;
      stage_57_active <= stage_56_active;
      stage_57_at_iter_0 <= stage_56_at_iter_0;
      stage_58_active <= stage_57_active;
      stage_58_at_iter_0 <= stage_57_at_iter_0;
      stage_59_active <= stage_58_active;
      stage_59_at_iter_0 <= stage_58_at_iter_0;
      stage_60_active <= stage_59_active;
      stage_60_at_iter_0 <= stage_59_at_iter_0;
      stage_61_active <= stage_60_active;
      stage_61_at_iter_0 <= stage_60_at_iter_0;
      stage_62_active <= stage_61_active;
      stage_62_at_iter_0 <= stage_61_at_iter_0;
      stage_63_active <= stage_62_active;
      stage_63_at_iter_0 <= stage_62_at_iter_0;
      stage_64_active <= stage_63_active;
      stage_64_at_iter_0 <= stage_63_at_iter_0;
      stage_65_active <= stage_64_active;
      stage_65_at_iter_0 <= stage_64_at_iter_0;
      stage_66_active <= stage_65_active;
      stage_66_at_iter_0 <= stage_65_at_iter_0;
      stage_67_active <= stage_66_active;
      stage_67_at_iter_0 <= stage_66_at_iter_0;
      stage_68_active <= stage_67_active;
      stage_68_at_iter_0 <= stage_67_at_iter_0;
      stage_69_active <= stage_68_active;
      stage_69_at_iter_0 <= stage_68_at_iter_0;
      stage_70_active <= stage_69_active;
      stage_70_at_iter_0 <= stage_69_at_iter_0;
      stage_71_active <= stage_70_active;
      stage_71_at_iter_0 <= stage_70_at_iter_0;
      stage_72_active <= stage_71_active;
      stage_72_at_iter_0 <= stage_71_at_iter_0;
      stage_73_active <= stage_72_active;
      stage_73_at_iter_0 <= stage_72_at_iter_0;
      stage_74_active <= stage_73_active;
      stage_74_at_iter_0 <= stage_73_at_iter_0;
      stage_75_active <= stage_74_active;
      stage_75_at_iter_0 <= stage_74_at_iter_0;
      stage_76_active <= stage_75_active;
      stage_76_at_iter_0 <= stage_75_at_iter_0;
      stage_77_active <= stage_76_active;
      stage_77_at_iter_0 <= stage_76_at_iter_0;
      stage_78_active <= stage_77_active;
      stage_78_at_iter_0 <= stage_77_at_iter_0;
      stage_79_active <= stage_78_active;
      stage_79_at_iter_0 <= stage_78_at_iter_0;
      stage_80_active <= stage_79_active;
      stage_80_at_iter_0 <= stage_79_at_iter_0;
      stage_81_active <= stage_80_active;
      stage_81_at_iter_0 <= stage_80_at_iter_0;
      stage_82_active <= stage_81_active;
      stage_82_at_iter_0 <= stage_81_at_iter_0;
      stage_83_active <= stage_82_active;
      stage_83_at_iter_0 <= stage_82_at_iter_0;
      stage_84_active <= stage_83_active;
      stage_84_at_iter_0 <= stage_83_at_iter_0;
      stage_85_active <= stage_84_active;
      stage_85_at_iter_0 <= stage_84_at_iter_0;
      stage_86_active <= stage_85_active;
      stage_86_at_iter_0 <= stage_85_at_iter_0;
      stage_87_active <= stage_86_active;
      stage_87_at_iter_0 <= stage_86_at_iter_0;
      stage_88_active <= stage_87_active;
      stage_88_at_iter_0 <= stage_87_at_iter_0;
      stage_89_active <= stage_88_active;
      stage_89_at_iter_0 <= stage_88_at_iter_0;
      stage_90_active <= stage_89_active;
      stage_90_at_iter_0 <= stage_89_at_iter_0;
      stage_91_active <= stage_90_active;
      stage_91_at_iter_0 <= stage_90_at_iter_0;
      stage_92_active <= stage_91_active;
      stage_92_at_iter_0 <= stage_91_at_iter_0;
      stage_93_active <= stage_92_active;
      stage_93_at_iter_0 <= stage_92_at_iter_0;
      stage_94_active <= stage_93_active;
      stage_94_at_iter_0 <= stage_93_at_iter_0;
      stage_95_active <= stage_94_active;
      stage_95_at_iter_0 <= stage_94_at_iter_0;
      stage_96_active <= stage_95_active;
      stage_96_at_iter_0 <= stage_95_at_iter_0;
      stage_97_active <= stage_96_active;
      stage_97_at_iter_0 <= stage_96_at_iter_0;
      stage_98_active <= stage_97_active;
      stage_98_at_iter_0 <= stage_97_at_iter_0;
      stage_99_active <= stage_98_active;
      stage_99_at_iter_0 <= stage_98_at_iter_0;
      stage_100_active <= stage_99_active;
      stage_100_at_iter_0 <= stage_99_at_iter_0;
      stage_101_active <= stage_100_active;
      stage_101_at_iter_0 <= stage_100_at_iter_0;
      stage_102_active <= stage_101_active;
      stage_102_at_iter_0 <= stage_101_at_iter_0;
      stage_103_active <= stage_102_active;
      stage_103_at_iter_0 <= stage_102_at_iter_0;
      stage_104_active <= stage_103_active;
      stage_104_at_iter_0 <= stage_103_at_iter_0;
      stage_105_active <= stage_104_active;
      stage_105_at_iter_0 <= stage_104_at_iter_0;
      stage_106_active <= stage_105_active;
      stage_106_at_iter_0 <= stage_105_at_iter_0;
      stage_107_active <= stage_106_active;
      stage_107_at_iter_0 <= stage_106_at_iter_0;
      stage_108_active <= stage_107_active;
      stage_108_at_iter_0 <= stage_107_at_iter_0;
      stage_109_active <= stage_108_active;
      stage_109_at_iter_0 <= stage_108_at_iter_0;
      stage_110_active <= stage_109_active;
      stage_110_at_iter_0 <= stage_109_at_iter_0;
      stage_111_active <= stage_110_active;
      stage_111_at_iter_0 <= stage_110_at_iter_0;
      stage_112_active <= stage_111_active;
      stage_112_at_iter_0 <= stage_111_at_iter_0;
      stage_113_active <= stage_112_active;
      stage_113_at_iter_0 <= stage_112_at_iter_0;
      stage_114_active <= stage_113_active;
      stage_114_at_iter_0 <= stage_113_at_iter_0;
      stage_115_active <= stage_114_active;
      stage_115_at_iter_0 <= stage_114_at_iter_0;
      stage_116_active <= stage_115_active;
      stage_116_at_iter_0 <= stage_115_at_iter_0;
      stage_117_active <= stage_116_active;
      stage_117_at_iter_0 <= stage_116_at_iter_0;
      stage_118_active <= stage_117_active;
      stage_118_at_iter_0 <= stage_117_at_iter_0;
      stage_119_active <= stage_118_active;
      stage_119_at_iter_0 <= stage_118_at_iter_0;
      stage_120_active <= stage_119_active;
      stage_120_at_iter_0 <= stage_119_at_iter_0;
      stage_121_active <= stage_120_active;
      stage_121_at_iter_0 <= stage_120_at_iter_0;
      stage_122_active <= stage_121_active;
      stage_122_at_iter_0 <= stage_121_at_iter_0;
      stage_123_active <= stage_122_active;
      stage_123_at_iter_0 <= stage_122_at_iter_0;
      stage_124_active <= stage_123_active;
      stage_124_at_iter_0 <= stage_123_at_iter_0;
      stage_125_active <= stage_124_active;
      stage_125_at_iter_0 <= stage_124_at_iter_0;
      stage_126_active <= stage_125_active;
      stage_126_at_iter_0 <= stage_125_at_iter_0;
      stage_127_active <= stage_126_active;
      stage_127_at_iter_0 <= stage_126_at_iter_0;
      stage_128_active <= stage_127_active;
      stage_128_at_iter_0 <= stage_127_at_iter_0;
      stage_129_active <= stage_128_active;
      stage_129_at_iter_0 <= stage_128_at_iter_0;
      stage_130_active <= stage_129_active;
      stage_130_at_iter_0 <= stage_129_at_iter_0;
      stage_131_active <= stage_130_active;
      stage_131_at_iter_0 <= stage_130_at_iter_0;
      stage_132_active <= stage_131_active;
      stage_132_at_iter_0 <= stage_131_at_iter_0;
      stage_133_active <= stage_132_active;
      stage_133_at_iter_0 <= stage_132_at_iter_0;
      stage_134_active <= stage_133_active;
      stage_134_at_iter_0 <= stage_133_at_iter_0;
      stage_135_active <= stage_134_active;
      stage_135_at_iter_0 <= stage_134_at_iter_0;
      stage_136_active <= stage_135_active;
      stage_136_at_iter_0 <= stage_135_at_iter_0;
      stage_137_active <= stage_136_active;
      stage_137_at_iter_0 <= stage_136_at_iter_0;
      stage_138_active <= stage_137_active;
      stage_138_at_iter_0 <= stage_137_at_iter_0;
      stage_139_active <= stage_138_active;
      stage_139_at_iter_0 <= stage_138_at_iter_0;
      stage_140_active <= stage_139_active;
      stage_140_at_iter_0 <= stage_139_at_iter_0;
      stage_141_active <= stage_140_active;
      stage_141_at_iter_0 <= stage_140_at_iter_0;
      stage_142_active <= stage_141_active;
      stage_142_at_iter_0 <= stage_141_at_iter_0;
      stage_143_active <= stage_142_active;
      stage_143_at_iter_0 <= stage_142_at_iter_0;
      stage_144_active <= stage_143_active;
      stage_144_at_iter_0 <= stage_143_at_iter_0;
      stage_145_active <= stage_144_active;
      stage_145_at_iter_0 <= stage_144_at_iter_0;
      stage_146_active <= stage_145_active;
      stage_146_at_iter_0 <= stage_145_at_iter_0;
      stage_147_active <= stage_146_active;
      stage_147_at_iter_0 <= stage_146_at_iter_0;
      stage_148_active <= stage_147_active;
      stage_148_at_iter_0 <= stage_147_at_iter_0;
      stage_149_active <= stage_148_active;
      stage_149_at_iter_0 <= stage_148_at_iter_0;
      stage_150_active <= stage_149_active;
      stage_150_at_iter_0 <= stage_149_at_iter_0;
      stage_151_active <= stage_150_active;
      stage_151_at_iter_0 <= stage_150_at_iter_0;
      stage_152_active <= stage_151_active;
      stage_152_at_iter_0 <= stage_151_at_iter_0;
      stage_153_active <= stage_152_active;
      stage_153_at_iter_0 <= stage_152_at_iter_0;
      stage_154_active <= stage_153_active;
      stage_154_at_iter_0 <= stage_153_at_iter_0;
      stage_155_active <= stage_154_active;
      stage_155_at_iter_0 <= stage_154_at_iter_0;
      stage_156_active <= stage_155_active;
      stage_156_at_iter_0 <= stage_155_at_iter_0;
      stage_157_active <= stage_156_active;
      stage_157_at_iter_0 <= stage_156_at_iter_0;
      stage_158_active <= stage_157_active;
      stage_158_at_iter_0 <= stage_157_at_iter_0;
      stage_159_active <= stage_158_active;
      stage_159_at_iter_0 <= stage_158_at_iter_0;
      stage_160_active <= stage_159_active;
      stage_160_at_iter_0 <= stage_159_at_iter_0;
      stage_161_active <= stage_160_active;
      stage_161_at_iter_0 <= stage_160_at_iter_0;
      stage_162_active <= stage_161_active;
      stage_162_at_iter_0 <= stage_161_at_iter_0;
      stage_163_active <= stage_162_active;
      stage_163_at_iter_0 <= stage_162_at_iter_0;
      stage_164_active <= stage_163_active;
      stage_164_at_iter_0 <= stage_163_at_iter_0;
      stage_165_active <= stage_164_active;
      stage_165_at_iter_0 <= stage_164_at_iter_0;
      stage_166_active <= stage_165_active;
      stage_166_at_iter_0 <= stage_165_at_iter_0;
      stage_167_active <= stage_166_active;
      stage_167_at_iter_0 <= stage_166_at_iter_0;
      stage_168_active <= stage_167_active;
      stage_168_at_iter_0 <= stage_167_at_iter_0;
      stage_169_active <= stage_168_active;
      stage_169_at_iter_0 <= stage_168_at_iter_0;
      stage_170_active <= stage_169_active;
      stage_170_at_iter_0 <= stage_169_at_iter_0;
      stage_171_active <= stage_170_active;
      stage_171_at_iter_0 <= stage_170_at_iter_0;
      stage_172_active <= stage_171_active;
      stage_172_at_iter_0 <= stage_171_at_iter_0;
      stage_173_active <= stage_172_active;
      stage_173_at_iter_0 <= stage_172_at_iter_0;
      stage_174_active <= stage_173_active;
      stage_174_at_iter_0 <= stage_173_at_iter_0;
      stage_175_active <= stage_174_active;
      stage_175_at_iter_0 <= stage_174_at_iter_0;
      stage_176_active <= stage_175_active;
      stage_176_at_iter_0 <= stage_175_at_iter_0;
      stage_177_active <= stage_176_active;
      stage_177_at_iter_0 <= stage_176_at_iter_0;
      stage_178_active <= stage_177_active;
      stage_178_at_iter_0 <= stage_177_at_iter_0;
      stage_179_active <= stage_178_active;
      stage_179_at_iter_0 <= stage_178_at_iter_0;
      stage_180_active <= stage_179_active;
      stage_180_at_iter_0 <= stage_179_at_iter_0;

      in_off_chip_in_update_0_read_read_0_stage_2 <= in_off_chip_in_update_0_read_read_0;
      in_off_chip_in_update_0_read_read_0_stage_3 <= in_off_chip_in_update_0_read_read_0_stage_2;
      in_off_chip_in_update_0_read_read_0_stage_4 <= in_off_chip_in_update_0_read_read_0_stage_3;
      in_off_chip_in_update_0_read_read_0_stage_5 <= in_off_chip_in_update_0_read_read_0_stage_4;
      in_off_chip_in_update_0_read_read_0_stage_6 <= in_off_chip_in_update_0_read_read_0_stage_5;
      in_off_chip_in_update_0_read_read_0_stage_7 <= in_off_chip_in_update_0_read_read_0_stage_6;
      in_off_chip_in_update_0_read_read_0_stage_8 <= in_off_chip_in_update_0_read_read_0_stage_7;
      in_off_chip_in_update_0_read_read_0_stage_9 <= in_off_chip_in_update_0_read_read_0_stage_8;
      in_off_chip_in_update_0_read_read_0_stage_10 <= in_off_chip_in_update_0_read_read_0_stage_9;
      in_off_chip_in_update_0_read_read_0_stage_11 <= in_off_chip_in_update_0_read_read_0_stage_10;
      in_off_chip_in_update_0_read_read_0_stage_12 <= in_off_chip_in_update_0_read_read_0_stage_11;
      in_off_chip_in_update_0_read_read_0_stage_13 <= in_off_chip_in_update_0_read_read_0_stage_12;
      in_off_chip_in_update_0_read_read_0_stage_14 <= in_off_chip_in_update_0_read_read_0_stage_13;
      in_off_chip_in_update_0_read_read_0_stage_15 <= in_off_chip_in_update_0_read_read_0_stage_14;
      in_off_chip_in_update_0_read_read_0_stage_16 <= in_off_chip_in_update_0_read_read_0_stage_15;
      in_off_chip_in_update_0_read_read_0_stage_17 <= in_off_chip_in_update_0_read_read_0_stage_16;
      in_off_chip_in_update_0_read_read_0_stage_18 <= in_off_chip_in_update_0_read_read_0_stage_17;
      in_off_chip_in_update_0_read_read_0_stage_19 <= in_off_chip_in_update_0_read_read_0_stage_18;
      in_off_chip_in_update_0_read_read_0_stage_20 <= in_off_chip_in_update_0_read_read_0_stage_19;
      in_off_chip_in_update_0_read_read_0_stage_21 <= in_off_chip_in_update_0_read_read_0_stage_20;
      in_off_chip_in_update_0_read_read_0_stage_22 <= in_off_chip_in_update_0_read_read_0_stage_21;
      in_off_chip_in_update_0_read_read_0_stage_23 <= in_off_chip_in_update_0_read_read_0_stage_22;
      in_off_chip_in_update_0_read_read_0_stage_24 <= in_off_chip_in_update_0_read_read_0_stage_23;
      in_off_chip_in_update_0_read_read_0_stage_25 <= in_off_chip_in_update_0_read_read_0_stage_24;
      in_off_chip_in_update_0_read_read_0_stage_26 <= in_off_chip_in_update_0_read_read_0_stage_25;
      in_off_chip_in_update_0_read_read_0_stage_27 <= in_off_chip_in_update_0_read_read_0_stage_26;
      in_off_chip_in_update_0_read_read_0_stage_28 <= in_off_chip_in_update_0_read_read_0_stage_27;
      in_off_chip_in_update_0_read_read_0_stage_29 <= in_off_chip_in_update_0_read_read_0_stage_28;
      in_off_chip_in_update_0_read_read_0_stage_30 <= in_off_chip_in_update_0_read_read_0_stage_29;
      in_off_chip_in_update_0_read_read_0_stage_31 <= in_off_chip_in_update_0_read_read_0_stage_30;
      in_off_chip_in_update_0_read_read_0_stage_32 <= in_off_chip_in_update_0_read_read_0_stage_31;
      in_off_chip_in_update_0_read_read_0_stage_33 <= in_off_chip_in_update_0_read_read_0_stage_32;
      in_off_chip_in_update_0_read_read_0_stage_34 <= in_off_chip_in_update_0_read_read_0_stage_33;
      in_off_chip_in_update_0_read_read_0_stage_35 <= in_off_chip_in_update_0_read_read_0_stage_34;
      in_off_chip_in_update_0_read_read_0_stage_36 <= in_off_chip_in_update_0_read_read_0_stage_35;
      in_off_chip_in_update_0_read_read_0_stage_37 <= in_off_chip_in_update_0_read_read_0_stage_36;
      in_off_chip_in_update_0_read_read_0_stage_38 <= in_off_chip_in_update_0_read_read_0_stage_37;
      in_off_chip_in_update_0_read_read_0_stage_39 <= in_off_chip_in_update_0_read_read_0_stage_38;
      in_off_chip_in_update_0_read_read_0_stage_40 <= in_off_chip_in_update_0_read_read_0_stage_39;
      in_off_chip_in_update_0_read_read_0_stage_41 <= in_off_chip_in_update_0_read_read_0_stage_40;
      in_off_chip_in_update_0_read_read_0_stage_42 <= in_off_chip_in_update_0_read_read_0_stage_41;
      in_off_chip_in_update_0_read_read_0_stage_43 <= in_off_chip_in_update_0_read_read_0_stage_42;
      in_off_chip_in_update_0_read_read_0_stage_44 <= in_off_chip_in_update_0_read_read_0_stage_43;
      in_off_chip_in_update_0_read_read_0_stage_45 <= in_off_chip_in_update_0_read_read_0_stage_44;
      in_off_chip_in_update_0_read_read_0_stage_46 <= in_off_chip_in_update_0_read_read_0_stage_45;
      in_off_chip_in_update_0_read_read_0_stage_47 <= in_off_chip_in_update_0_read_read_0_stage_46;
      in_off_chip_in_update_0_read_read_0_stage_48 <= in_off_chip_in_update_0_read_read_0_stage_47;
      in_off_chip_in_update_0_read_read_0_stage_49 <= in_off_chip_in_update_0_read_read_0_stage_48;
      in_off_chip_in_update_0_read_read_0_stage_50 <= in_off_chip_in_update_0_read_read_0_stage_49;
      in_off_chip_in_update_0_read_read_0_stage_51 <= in_off_chip_in_update_0_read_read_0_stage_50;
      in_off_chip_in_update_0_read_read_0_stage_52 <= in_off_chip_in_update_0_read_read_0_stage_51;
      in_off_chip_in_update_0_read_read_0_stage_53 <= in_off_chip_in_update_0_read_read_0_stage_52;
      in_off_chip_in_update_0_read_read_0_stage_54 <= in_off_chip_in_update_0_read_read_0_stage_53;
      in_off_chip_in_update_0_read_read_0_stage_55 <= in_off_chip_in_update_0_read_read_0_stage_54;
      in_off_chip_in_update_0_read_read_0_stage_56 <= in_off_chip_in_update_0_read_read_0_stage_55;
      in_off_chip_in_update_0_read_read_0_stage_57 <= in_off_chip_in_update_0_read_read_0_stage_56;
      in_off_chip_in_update_0_read_read_0_stage_58 <= in_off_chip_in_update_0_read_read_0_stage_57;
      in_off_chip_in_update_0_read_read_0_stage_59 <= in_off_chip_in_update_0_read_read_0_stage_58;
      in_off_chip_in_update_0_read_read_0_stage_60 <= in_off_chip_in_update_0_read_read_0_stage_59;
      in_off_chip_in_update_0_read_read_0_stage_61 <= in_off_chip_in_update_0_read_read_0_stage_60;
      in_off_chip_in_update_0_read_read_0_stage_62 <= in_off_chip_in_update_0_read_read_0_stage_61;
      in_off_chip_in_update_0_read_read_0_stage_63 <= in_off_chip_in_update_0_read_read_0_stage_62;
      in_off_chip_in_update_0_read_read_0_stage_64 <= in_off_chip_in_update_0_read_read_0_stage_63;
      in_off_chip_in_update_0_read_read_0_stage_65 <= in_off_chip_in_update_0_read_read_0_stage_64;
      in_off_chip_in_update_0_read_read_0_stage_66 <= in_off_chip_in_update_0_read_read_0_stage_65;
      in_off_chip_in_update_0_read_read_0_stage_67 <= in_off_chip_in_update_0_read_read_0_stage_66;
      in_off_chip_in_update_0_read_read_0_stage_68 <= in_off_chip_in_update_0_read_read_0_stage_67;
      in_off_chip_in_update_0_read_read_0_stage_69 <= in_off_chip_in_update_0_read_read_0_stage_68;
      in_off_chip_in_update_0_read_read_0_stage_70 <= in_off_chip_in_update_0_read_read_0_stage_69;
      in_off_chip_in_update_0_read_read_0_stage_71 <= in_off_chip_in_update_0_read_read_0_stage_70;
      in_off_chip_in_update_0_read_read_0_stage_72 <= in_off_chip_in_update_0_read_read_0_stage_71;
      in_off_chip_in_update_0_read_read_0_stage_73 <= in_off_chip_in_update_0_read_read_0_stage_72;
      in_off_chip_in_update_0_read_read_0_stage_74 <= in_off_chip_in_update_0_read_read_0_stage_73;
      in_off_chip_in_update_0_read_read_0_stage_75 <= in_off_chip_in_update_0_read_read_0_stage_74;
      in_off_chip_in_update_0_read_read_0_stage_76 <= in_off_chip_in_update_0_read_read_0_stage_75;
      in_off_chip_in_update_0_read_read_0_stage_77 <= in_off_chip_in_update_0_read_read_0_stage_76;
      in_off_chip_in_update_0_read_read_0_stage_78 <= in_off_chip_in_update_0_read_read_0_stage_77;
      in_off_chip_in_update_0_read_read_0_stage_79 <= in_off_chip_in_update_0_read_read_0_stage_78;
      in_off_chip_in_update_0_read_read_0_stage_80 <= in_off_chip_in_update_0_read_read_0_stage_79;
      in_off_chip_in_update_0_read_read_0_stage_81 <= in_off_chip_in_update_0_read_read_0_stage_80;
      in_off_chip_in_update_0_read_read_0_stage_82 <= in_off_chip_in_update_0_read_read_0_stage_81;
      in_off_chip_in_update_0_read_read_0_stage_83 <= in_off_chip_in_update_0_read_read_0_stage_82;
      in_off_chip_in_update_0_read_read_0_stage_84 <= in_off_chip_in_update_0_read_read_0_stage_83;
      in_off_chip_in_update_0_read_read_0_stage_85 <= in_off_chip_in_update_0_read_read_0_stage_84;
      in_off_chip_in_update_0_read_read_0_stage_86 <= in_off_chip_in_update_0_read_read_0_stage_85;
      in_off_chip_in_update_0_read_read_0_stage_87 <= in_off_chip_in_update_0_read_read_0_stage_86;
      in_off_chip_in_update_0_read_read_0_stage_88 <= in_off_chip_in_update_0_read_read_0_stage_87;
      in_off_chip_in_update_0_read_read_0_stage_89 <= in_off_chip_in_update_0_read_read_0_stage_88;
      in_off_chip_in_update_0_read_read_0_stage_90 <= in_off_chip_in_update_0_read_read_0_stage_89;
      in_off_chip_in_update_0_read_read_0_stage_91 <= in_off_chip_in_update_0_read_read_0_stage_90;
      in_off_chip_in_update_0_read_read_0_stage_92 <= in_off_chip_in_update_0_read_read_0_stage_91;
      in_off_chip_in_update_0_read_read_0_stage_93 <= in_off_chip_in_update_0_read_read_0_stage_92;
      in_off_chip_in_update_0_read_read_0_stage_94 <= in_off_chip_in_update_0_read_read_0_stage_93;
      in_off_chip_in_update_0_read_read_0_stage_95 <= in_off_chip_in_update_0_read_read_0_stage_94;
      in_off_chip_in_update_0_read_read_0_stage_96 <= in_off_chip_in_update_0_read_read_0_stage_95;
      in_off_chip_in_update_0_read_read_0_stage_97 <= in_off_chip_in_update_0_read_read_0_stage_96;
      in_off_chip_in_update_0_read_read_0_stage_98 <= in_off_chip_in_update_0_read_read_0_stage_97;
      in_off_chip_in_update_0_read_read_0_stage_99 <= in_off_chip_in_update_0_read_read_0_stage_98;
      in_off_chip_in_update_0_read_read_0_stage_100 <= in_off_chip_in_update_0_read_read_0_stage_99;
      in_off_chip_in_update_0_read_read_0_stage_101 <= in_off_chip_in_update_0_read_read_0_stage_100;
      in_off_chip_in_update_0_read_read_0_stage_102 <= in_off_chip_in_update_0_read_read_0_stage_101;
      in_off_chip_in_update_0_read_read_0_stage_103 <= in_off_chip_in_update_0_read_read_0_stage_102;
      in_off_chip_in_update_0_read_read_0_stage_104 <= in_off_chip_in_update_0_read_read_0_stage_103;
      in_off_chip_in_update_0_read_read_0_stage_105 <= in_off_chip_in_update_0_read_read_0_stage_104;
      in_off_chip_in_update_0_read_read_0_stage_106 <= in_off_chip_in_update_0_read_read_0_stage_105;
      in_off_chip_in_update_0_read_read_0_stage_107 <= in_off_chip_in_update_0_read_read_0_stage_106;
      in_off_chip_in_update_0_read_read_0_stage_108 <= in_off_chip_in_update_0_read_read_0_stage_107;
      in_off_chip_in_update_0_read_read_0_stage_109 <= in_off_chip_in_update_0_read_read_0_stage_108;
      in_off_chip_in_update_0_read_read_0_stage_110 <= in_off_chip_in_update_0_read_read_0_stage_109;
      in_off_chip_in_update_0_read_read_0_stage_111 <= in_off_chip_in_update_0_read_read_0_stage_110;
      in_off_chip_in_update_0_read_read_0_stage_112 <= in_off_chip_in_update_0_read_read_0_stage_111;
      in_off_chip_in_update_0_read_read_0_stage_113 <= in_off_chip_in_update_0_read_read_0_stage_112;
      in_off_chip_in_update_0_read_read_0_stage_114 <= in_off_chip_in_update_0_read_read_0_stage_113;
      in_off_chip_in_update_0_read_read_0_stage_115 <= in_off_chip_in_update_0_read_read_0_stage_114;
      in_off_chip_in_update_0_read_read_0_stage_116 <= in_off_chip_in_update_0_read_read_0_stage_115;
      in_off_chip_in_update_0_read_read_0_stage_117 <= in_off_chip_in_update_0_read_read_0_stage_116;
      in_off_chip_in_update_0_read_read_0_stage_118 <= in_off_chip_in_update_0_read_read_0_stage_117;
      in_off_chip_in_update_0_read_read_0_stage_119 <= in_off_chip_in_update_0_read_read_0_stage_118;
      in_off_chip_in_update_0_read_read_0_stage_120 <= in_off_chip_in_update_0_read_read_0_stage_119;
      in_off_chip_in_update_0_read_read_0_stage_121 <= in_off_chip_in_update_0_read_read_0_stage_120;
      in_off_chip_in_update_0_read_read_0_stage_122 <= in_off_chip_in_update_0_read_read_0_stage_121;
      in_off_chip_in_update_0_read_read_0_stage_123 <= in_off_chip_in_update_0_read_read_0_stage_122;
      in_off_chip_in_update_0_read_read_0_stage_124 <= in_off_chip_in_update_0_read_read_0_stage_123;
      in_off_chip_in_update_0_read_read_0_stage_125 <= in_off_chip_in_update_0_read_read_0_stage_124;
      in_off_chip_in_update_0_read_read_0_stage_126 <= in_off_chip_in_update_0_read_read_0_stage_125;
      in_off_chip_in_update_0_read_read_0_stage_127 <= in_off_chip_in_update_0_read_read_0_stage_126;
      in_off_chip_in_update_0_read_read_0_stage_128 <= in_off_chip_in_update_0_read_read_0_stage_127;
      in_off_chip_in_update_0_read_read_0_stage_129 <= in_off_chip_in_update_0_read_read_0_stage_128;
      in_off_chip_in_update_0_read_read_0_stage_130 <= in_off_chip_in_update_0_read_read_0_stage_129;
      in_off_chip_in_update_0_read_read_0_stage_131 <= in_off_chip_in_update_0_read_read_0_stage_130;
      in_off_chip_in_update_0_read_read_0_stage_132 <= in_off_chip_in_update_0_read_read_0_stage_131;
      in_off_chip_in_update_0_read_read_0_stage_133 <= in_off_chip_in_update_0_read_read_0_stage_132;
      in_off_chip_in_update_0_read_read_0_stage_134 <= in_off_chip_in_update_0_read_read_0_stage_133;
      in_off_chip_in_update_0_read_read_0_stage_135 <= in_off_chip_in_update_0_read_read_0_stage_134;
      in_off_chip_in_update_0_read_read_0_stage_136 <= in_off_chip_in_update_0_read_read_0_stage_135;
      in_off_chip_in_update_0_read_read_0_stage_137 <= in_off_chip_in_update_0_read_read_0_stage_136;
      in_off_chip_in_update_0_read_read_0_stage_138 <= in_off_chip_in_update_0_read_read_0_stage_137;
      in_off_chip_in_update_0_read_read_0_stage_139 <= in_off_chip_in_update_0_read_read_0_stage_138;
      in_off_chip_in_update_0_read_read_0_stage_140 <= in_off_chip_in_update_0_read_read_0_stage_139;
      in_off_chip_in_update_0_read_read_0_stage_141 <= in_off_chip_in_update_0_read_read_0_stage_140;
      in_off_chip_in_update_0_read_read_0_stage_142 <= in_off_chip_in_update_0_read_read_0_stage_141;
      in_off_chip_in_update_0_read_read_0_stage_143 <= in_off_chip_in_update_0_read_read_0_stage_142;
      in_off_chip_in_update_0_read_read_0_stage_144 <= in_off_chip_in_update_0_read_read_0_stage_143;
      in_off_chip_in_update_0_read_read_0_stage_145 <= in_off_chip_in_update_0_read_read_0_stage_144;
      in_off_chip_in_update_0_read_read_0_stage_146 <= in_off_chip_in_update_0_read_read_0_stage_145;
      in_off_chip_in_update_0_read_read_0_stage_147 <= in_off_chip_in_update_0_read_read_0_stage_146;
      in_off_chip_in_update_0_read_read_0_stage_148 <= in_off_chip_in_update_0_read_read_0_stage_147;
      in_off_chip_in_update_0_read_read_0_stage_149 <= in_off_chip_in_update_0_read_read_0_stage_148;
      in_off_chip_in_update_0_read_read_0_stage_150 <= in_off_chip_in_update_0_read_read_0_stage_149;
      in_off_chip_in_update_0_read_read_0_stage_151 <= in_off_chip_in_update_0_read_read_0_stage_150;
      in_off_chip_in_update_0_read_read_0_stage_152 <= in_off_chip_in_update_0_read_read_0_stage_151;
      in_off_chip_in_update_0_read_read_0_stage_153 <= in_off_chip_in_update_0_read_read_0_stage_152;
      in_off_chip_in_update_0_read_read_0_stage_154 <= in_off_chip_in_update_0_read_read_0_stage_153;
      in_off_chip_in_update_0_read_read_0_stage_155 <= in_off_chip_in_update_0_read_read_0_stage_154;
      in_off_chip_in_update_0_read_read_0_stage_156 <= in_off_chip_in_update_0_read_read_0_stage_155;
      in_off_chip_in_update_0_read_read_0_stage_157 <= in_off_chip_in_update_0_read_read_0_stage_156;
      in_off_chip_in_update_0_read_read_0_stage_158 <= in_off_chip_in_update_0_read_read_0_stage_157;
      in_off_chip_in_update_0_read_read_0_stage_159 <= in_off_chip_in_update_0_read_read_0_stage_158;
      in_off_chip_in_update_0_read_read_0_stage_160 <= in_off_chip_in_update_0_read_read_0_stage_159;
      in_off_chip_in_update_0_read_read_0_stage_161 <= in_off_chip_in_update_0_read_read_0_stage_160;
      in_off_chip_in_update_0_read_read_0_stage_162 <= in_off_chip_in_update_0_read_read_0_stage_161;
      in_off_chip_in_update_0_read_read_0_stage_163 <= in_off_chip_in_update_0_read_read_0_stage_162;
      in_off_chip_in_update_0_read_read_0_stage_164 <= in_off_chip_in_update_0_read_read_0_stage_163;
      in_off_chip_in_update_0_read_read_0_stage_165 <= in_off_chip_in_update_0_read_read_0_stage_164;
      in_off_chip_in_update_0_read_read_0_stage_166 <= in_off_chip_in_update_0_read_read_0_stage_165;
      in_off_chip_in_update_0_read_read_0_stage_167 <= in_off_chip_in_update_0_read_read_0_stage_166;
      in_off_chip_in_update_0_read_read_0_stage_168 <= in_off_chip_in_update_0_read_read_0_stage_167;
      in_off_chip_in_update_0_read_read_0_stage_169 <= in_off_chip_in_update_0_read_read_0_stage_168;
      in_off_chip_in_update_0_read_read_0_stage_170 <= in_off_chip_in_update_0_read_read_0_stage_169;
      in_off_chip_in_update_0_read_read_0_stage_171 <= in_off_chip_in_update_0_read_read_0_stage_170;
      in_off_chip_in_update_0_read_read_0_stage_172 <= in_off_chip_in_update_0_read_read_0_stage_171;
      in_off_chip_in_update_0_read_read_0_stage_173 <= in_off_chip_in_update_0_read_read_0_stage_172;
      in_off_chip_in_update_0_read_read_0_stage_174 <= in_off_chip_in_update_0_read_read_0_stage_173;
      in_off_chip_in_update_0_read_read_0_stage_175 <= in_off_chip_in_update_0_read_read_0_stage_174;
      in_off_chip_in_update_0_read_read_0_stage_176 <= in_off_chip_in_update_0_read_read_0_stage_175;
      in_off_chip_in_update_0_read_read_0_stage_177 <= in_off_chip_in_update_0_read_read_0_stage_176;
      in_off_chip_in_update_0_read_read_0_stage_178 <= in_off_chip_in_update_0_read_read_0_stage_177;
      in_off_chip_in_update_0_read_read_0_stage_179 <= in_off_chip_in_update_0_read_read_0_stage_178;
      in_off_chip_in_update_0_read_read_0_stage_180 <= in_off_chip_in_update_0_read_read_0_stage_179;
      in_off_chip_in_update_0_read_read_0_stage_181 <= in_off_chip_in_update_0_read_read_0_stage_180;
      in_update_0_stage_3 <= in_update_0;
      in_update_0_stage_4 <= in_update_0_stage_3;
      in_update_0_stage_5 <= in_update_0_stage_4;
      in_update_0_stage_6 <= in_update_0_stage_5;
      in_update_0_stage_7 <= in_update_0_stage_6;
      in_update_0_stage_8 <= in_update_0_stage_7;
      in_update_0_stage_9 <= in_update_0_stage_8;
      in_update_0_stage_10 <= in_update_0_stage_9;
      in_update_0_stage_11 <= in_update_0_stage_10;
      in_update_0_stage_12 <= in_update_0_stage_11;
      in_update_0_stage_13 <= in_update_0_stage_12;
      in_update_0_stage_14 <= in_update_0_stage_13;
      in_update_0_stage_15 <= in_update_0_stage_14;
      in_update_0_stage_16 <= in_update_0_stage_15;
      in_update_0_stage_17 <= in_update_0_stage_16;
      in_update_0_stage_18 <= in_update_0_stage_17;
      in_update_0_stage_19 <= in_update_0_stage_18;
      in_update_0_stage_20 <= in_update_0_stage_19;
      in_update_0_stage_21 <= in_update_0_stage_20;
      in_update_0_stage_22 <= in_update_0_stage_21;
      in_update_0_stage_23 <= in_update_0_stage_22;
      in_update_0_stage_24 <= in_update_0_stage_23;
      in_update_0_stage_25 <= in_update_0_stage_24;
      in_update_0_stage_26 <= in_update_0_stage_25;
      in_update_0_stage_27 <= in_update_0_stage_26;
      in_update_0_stage_28 <= in_update_0_stage_27;
      in_update_0_stage_29 <= in_update_0_stage_28;
      in_update_0_stage_30 <= in_update_0_stage_29;
      in_update_0_stage_31 <= in_update_0_stage_30;
      in_update_0_stage_32 <= in_update_0_stage_31;
      in_update_0_stage_33 <= in_update_0_stage_32;
      in_update_0_stage_34 <= in_update_0_stage_33;
      in_update_0_stage_35 <= in_update_0_stage_34;
      in_update_0_stage_36 <= in_update_0_stage_35;
      in_update_0_stage_37 <= in_update_0_stage_36;
      in_update_0_stage_38 <= in_update_0_stage_37;
      in_update_0_stage_39 <= in_update_0_stage_38;
      in_update_0_stage_40 <= in_update_0_stage_39;
      in_update_0_stage_41 <= in_update_0_stage_40;
      in_update_0_stage_42 <= in_update_0_stage_41;
      in_update_0_stage_43 <= in_update_0_stage_42;
      in_update_0_stage_44 <= in_update_0_stage_43;
      in_update_0_stage_45 <= in_update_0_stage_44;
      in_update_0_stage_46 <= in_update_0_stage_45;
      in_update_0_stage_47 <= in_update_0_stage_46;
      in_update_0_stage_48 <= in_update_0_stage_47;
      in_update_0_stage_49 <= in_update_0_stage_48;
      in_update_0_stage_50 <= in_update_0_stage_49;
      in_update_0_stage_51 <= in_update_0_stage_50;
      in_update_0_stage_52 <= in_update_0_stage_51;
      in_update_0_stage_53 <= in_update_0_stage_52;
      in_update_0_stage_54 <= in_update_0_stage_53;
      in_update_0_stage_55 <= in_update_0_stage_54;
      in_update_0_stage_56 <= in_update_0_stage_55;
      in_update_0_stage_57 <= in_update_0_stage_56;
      in_update_0_stage_58 <= in_update_0_stage_57;
      in_update_0_stage_59 <= in_update_0_stage_58;
      in_update_0_stage_60 <= in_update_0_stage_59;
      in_update_0_stage_61 <= in_update_0_stage_60;
      in_update_0_stage_62 <= in_update_0_stage_61;
      in_update_0_stage_63 <= in_update_0_stage_62;
      in_update_0_stage_64 <= in_update_0_stage_63;
      in_update_0_stage_65 <= in_update_0_stage_64;
      in_update_0_stage_66 <= in_update_0_stage_65;
      in_update_0_stage_67 <= in_update_0_stage_66;
      in_update_0_stage_68 <= in_update_0_stage_67;
      in_update_0_stage_69 <= in_update_0_stage_68;
      in_update_0_stage_70 <= in_update_0_stage_69;
      in_update_0_stage_71 <= in_update_0_stage_70;
      in_update_0_stage_72 <= in_update_0_stage_71;
      in_update_0_stage_73 <= in_update_0_stage_72;
      in_update_0_stage_74 <= in_update_0_stage_73;
      in_update_0_stage_75 <= in_update_0_stage_74;
      in_update_0_stage_76 <= in_update_0_stage_75;
      in_update_0_stage_77 <= in_update_0_stage_76;
      in_update_0_stage_78 <= in_update_0_stage_77;
      in_update_0_stage_79 <= in_update_0_stage_78;
      in_update_0_stage_80 <= in_update_0_stage_79;
      in_update_0_stage_81 <= in_update_0_stage_80;
      in_update_0_stage_82 <= in_update_0_stage_81;
      in_update_0_stage_83 <= in_update_0_stage_82;
      in_update_0_stage_84 <= in_update_0_stage_83;
      in_update_0_stage_85 <= in_update_0_stage_84;
      in_update_0_stage_86 <= in_update_0_stage_85;
      in_update_0_stage_87 <= in_update_0_stage_86;
      in_update_0_stage_88 <= in_update_0_stage_87;
      in_update_0_stage_89 <= in_update_0_stage_88;
      in_update_0_stage_90 <= in_update_0_stage_89;
      in_update_0_stage_91 <= in_update_0_stage_90;
      in_update_0_stage_92 <= in_update_0_stage_91;
      in_update_0_stage_93 <= in_update_0_stage_92;
      in_update_0_stage_94 <= in_update_0_stage_93;
      in_update_0_stage_95 <= in_update_0_stage_94;
      in_update_0_stage_96 <= in_update_0_stage_95;
      in_update_0_stage_97 <= in_update_0_stage_96;
      in_update_0_stage_98 <= in_update_0_stage_97;
      in_update_0_stage_99 <= in_update_0_stage_98;
      in_update_0_stage_100 <= in_update_0_stage_99;
      in_update_0_stage_101 <= in_update_0_stage_100;
      in_update_0_stage_102 <= in_update_0_stage_101;
      in_update_0_stage_103 <= in_update_0_stage_102;
      in_update_0_stage_104 <= in_update_0_stage_103;
      in_update_0_stage_105 <= in_update_0_stage_104;
      in_update_0_stage_106 <= in_update_0_stage_105;
      in_update_0_stage_107 <= in_update_0_stage_106;
      in_update_0_stage_108 <= in_update_0_stage_107;
      in_update_0_stage_109 <= in_update_0_stage_108;
      in_update_0_stage_110 <= in_update_0_stage_109;
      in_update_0_stage_111 <= in_update_0_stage_110;
      in_update_0_stage_112 <= in_update_0_stage_111;
      in_update_0_stage_113 <= in_update_0_stage_112;
      in_update_0_stage_114 <= in_update_0_stage_113;
      in_update_0_stage_115 <= in_update_0_stage_114;
      in_update_0_stage_116 <= in_update_0_stage_115;
      in_update_0_stage_117 <= in_update_0_stage_116;
      in_update_0_stage_118 <= in_update_0_stage_117;
      in_update_0_stage_119 <= in_update_0_stage_118;
      in_update_0_stage_120 <= in_update_0_stage_119;
      in_update_0_stage_121 <= in_update_0_stage_120;
      in_update_0_stage_122 <= in_update_0_stage_121;
      in_update_0_stage_123 <= in_update_0_stage_122;
      in_update_0_stage_124 <= in_update_0_stage_123;
      in_update_0_stage_125 <= in_update_0_stage_124;
      in_update_0_stage_126 <= in_update_0_stage_125;
      in_update_0_stage_127 <= in_update_0_stage_126;
      in_update_0_stage_128 <= in_update_0_stage_127;
      in_update_0_stage_129 <= in_update_0_stage_128;
      in_update_0_stage_130 <= in_update_0_stage_129;
      in_update_0_stage_131 <= in_update_0_stage_130;
      in_update_0_stage_132 <= in_update_0_stage_131;
      in_update_0_stage_133 <= in_update_0_stage_132;
      in_update_0_stage_134 <= in_update_0_stage_133;
      in_update_0_stage_135 <= in_update_0_stage_134;
      in_update_0_stage_136 <= in_update_0_stage_135;
      in_update_0_stage_137 <= in_update_0_stage_136;
      in_update_0_stage_138 <= in_update_0_stage_137;
      in_update_0_stage_139 <= in_update_0_stage_138;
      in_update_0_stage_140 <= in_update_0_stage_139;
      in_update_0_stage_141 <= in_update_0_stage_140;
      in_update_0_stage_142 <= in_update_0_stage_141;
      in_update_0_stage_143 <= in_update_0_stage_142;
      in_update_0_stage_144 <= in_update_0_stage_143;
      in_update_0_stage_145 <= in_update_0_stage_144;
      in_update_0_stage_146 <= in_update_0_stage_145;
      in_update_0_stage_147 <= in_update_0_stage_146;
      in_update_0_stage_148 <= in_update_0_stage_147;
      in_update_0_stage_149 <= in_update_0_stage_148;
      in_update_0_stage_150 <= in_update_0_stage_149;
      in_update_0_stage_151 <= in_update_0_stage_150;
      in_update_0_stage_152 <= in_update_0_stage_151;
      in_update_0_stage_153 <= in_update_0_stage_152;
      in_update_0_stage_154 <= in_update_0_stage_153;
      in_update_0_stage_155 <= in_update_0_stage_154;
      in_update_0_stage_156 <= in_update_0_stage_155;
      in_update_0_stage_157 <= in_update_0_stage_156;
      in_update_0_stage_158 <= in_update_0_stage_157;
      in_update_0_stage_159 <= in_update_0_stage_158;
      in_update_0_stage_160 <= in_update_0_stage_159;
      in_update_0_stage_161 <= in_update_0_stage_160;
      in_update_0_stage_162 <= in_update_0_stage_161;
      in_update_0_stage_163 <= in_update_0_stage_162;
      in_update_0_stage_164 <= in_update_0_stage_163;
      in_update_0_stage_165 <= in_update_0_stage_164;
      in_update_0_stage_166 <= in_update_0_stage_165;
      in_update_0_stage_167 <= in_update_0_stage_166;
      in_update_0_stage_168 <= in_update_0_stage_167;
      in_update_0_stage_169 <= in_update_0_stage_168;
      in_update_0_stage_170 <= in_update_0_stage_169;
      in_update_0_stage_171 <= in_update_0_stage_170;
      in_update_0_stage_172 <= in_update_0_stage_171;
      in_update_0_stage_173 <= in_update_0_stage_172;
      in_update_0_stage_174 <= in_update_0_stage_173;
      in_update_0_stage_175 <= in_update_0_stage_174;
      in_update_0_stage_176 <= in_update_0_stage_175;
      in_update_0_stage_177 <= in_update_0_stage_176;
      in_update_0_stage_178 <= in_update_0_stage_177;
      in_update_0_stage_179 <= in_update_0_stage_178;
      in_update_0_stage_180 <= in_update_0_stage_179;
      in_update_0_stage_181 <= in_update_0_stage_180;
      bright_bright_weights_update_0_read_read_4_stage_8 <= bright_bright_weights_update_0_read_read_4;
      bright_bright_weights_update_0_read_read_4_stage_9 <= bright_bright_weights_update_0_read_read_4_stage_8;
      bright_bright_weights_update_0_read_read_4_stage_10 <= bright_bright_weights_update_0_read_read_4_stage_9;
      bright_bright_weights_update_0_read_read_4_stage_11 <= bright_bright_weights_update_0_read_read_4_stage_10;
      bright_bright_weights_update_0_read_read_4_stage_12 <= bright_bright_weights_update_0_read_read_4_stage_11;
      bright_bright_weights_update_0_read_read_4_stage_13 <= bright_bright_weights_update_0_read_read_4_stage_12;
      bright_bright_weights_update_0_read_read_4_stage_14 <= bright_bright_weights_update_0_read_read_4_stage_13;
      bright_bright_weights_update_0_read_read_4_stage_15 <= bright_bright_weights_update_0_read_read_4_stage_14;
      bright_bright_weights_update_0_read_read_4_stage_16 <= bright_bright_weights_update_0_read_read_4_stage_15;
      bright_bright_weights_update_0_read_read_4_stage_17 <= bright_bright_weights_update_0_read_read_4_stage_16;
      bright_bright_weights_update_0_read_read_4_stage_18 <= bright_bright_weights_update_0_read_read_4_stage_17;
      bright_bright_weights_update_0_read_read_4_stage_19 <= bright_bright_weights_update_0_read_read_4_stage_18;
      bright_bright_weights_update_0_read_read_4_stage_20 <= bright_bright_weights_update_0_read_read_4_stage_19;
      bright_bright_weights_update_0_read_read_4_stage_21 <= bright_bright_weights_update_0_read_read_4_stage_20;
      bright_bright_weights_update_0_read_read_4_stage_22 <= bright_bright_weights_update_0_read_read_4_stage_21;
      bright_bright_weights_update_0_read_read_4_stage_23 <= bright_bright_weights_update_0_read_read_4_stage_22;
      bright_bright_weights_update_0_read_read_4_stage_24 <= bright_bright_weights_update_0_read_read_4_stage_23;
      bright_bright_weights_update_0_read_read_4_stage_25 <= bright_bright_weights_update_0_read_read_4_stage_24;
      bright_bright_weights_update_0_read_read_4_stage_26 <= bright_bright_weights_update_0_read_read_4_stage_25;
      bright_bright_weights_update_0_read_read_4_stage_27 <= bright_bright_weights_update_0_read_read_4_stage_26;
      bright_bright_weights_update_0_read_read_4_stage_28 <= bright_bright_weights_update_0_read_read_4_stage_27;
      bright_bright_weights_update_0_read_read_4_stage_29 <= bright_bright_weights_update_0_read_read_4_stage_28;
      bright_bright_weights_update_0_read_read_4_stage_30 <= bright_bright_weights_update_0_read_read_4_stage_29;
      bright_bright_weights_update_0_read_read_4_stage_31 <= bright_bright_weights_update_0_read_read_4_stage_30;
      bright_bright_weights_update_0_read_read_4_stage_32 <= bright_bright_weights_update_0_read_read_4_stage_31;
      bright_bright_weights_update_0_read_read_4_stage_33 <= bright_bright_weights_update_0_read_read_4_stage_32;
      bright_bright_weights_update_0_read_read_4_stage_34 <= bright_bright_weights_update_0_read_read_4_stage_33;
      bright_bright_weights_update_0_read_read_4_stage_35 <= bright_bright_weights_update_0_read_read_4_stage_34;
      bright_bright_weights_update_0_read_read_4_stage_36 <= bright_bright_weights_update_0_read_read_4_stage_35;
      bright_bright_weights_update_0_read_read_4_stage_37 <= bright_bright_weights_update_0_read_read_4_stage_36;
      bright_bright_weights_update_0_read_read_4_stage_38 <= bright_bright_weights_update_0_read_read_4_stage_37;
      bright_bright_weights_update_0_read_read_4_stage_39 <= bright_bright_weights_update_0_read_read_4_stage_38;
      bright_bright_weights_update_0_read_read_4_stage_40 <= bright_bright_weights_update_0_read_read_4_stage_39;
      bright_bright_weights_update_0_read_read_4_stage_41 <= bright_bright_weights_update_0_read_read_4_stage_40;
      bright_bright_weights_update_0_read_read_4_stage_42 <= bright_bright_weights_update_0_read_read_4_stage_41;
      bright_bright_weights_update_0_read_read_4_stage_43 <= bright_bright_weights_update_0_read_read_4_stage_42;
      bright_bright_weights_update_0_read_read_4_stage_44 <= bright_bright_weights_update_0_read_read_4_stage_43;
      bright_bright_weights_update_0_read_read_4_stage_45 <= bright_bright_weights_update_0_read_read_4_stage_44;
      bright_bright_weights_update_0_read_read_4_stage_46 <= bright_bright_weights_update_0_read_read_4_stage_45;
      bright_bright_weights_update_0_read_read_4_stage_47 <= bright_bright_weights_update_0_read_read_4_stage_46;
      bright_bright_weights_update_0_read_read_4_stage_48 <= bright_bright_weights_update_0_read_read_4_stage_47;
      bright_bright_weights_update_0_read_read_4_stage_49 <= bright_bright_weights_update_0_read_read_4_stage_48;
      bright_bright_weights_update_0_read_read_4_stage_50 <= bright_bright_weights_update_0_read_read_4_stage_49;
      bright_bright_weights_update_0_read_read_4_stage_51 <= bright_bright_weights_update_0_read_read_4_stage_50;
      bright_bright_weights_update_0_read_read_4_stage_52 <= bright_bright_weights_update_0_read_read_4_stage_51;
      bright_bright_weights_update_0_read_read_4_stage_53 <= bright_bright_weights_update_0_read_read_4_stage_52;
      bright_bright_weights_update_0_read_read_4_stage_54 <= bright_bright_weights_update_0_read_read_4_stage_53;
      bright_bright_weights_update_0_read_read_4_stage_55 <= bright_bright_weights_update_0_read_read_4_stage_54;
      bright_bright_weights_update_0_read_read_4_stage_56 <= bright_bright_weights_update_0_read_read_4_stage_55;
      bright_bright_weights_update_0_read_read_4_stage_57 <= bright_bright_weights_update_0_read_read_4_stage_56;
      bright_bright_weights_update_0_read_read_4_stage_58 <= bright_bright_weights_update_0_read_read_4_stage_57;
      bright_bright_weights_update_0_read_read_4_stage_59 <= bright_bright_weights_update_0_read_read_4_stage_58;
      bright_bright_weights_update_0_read_read_4_stage_60 <= bright_bright_weights_update_0_read_read_4_stage_59;
      bright_bright_weights_update_0_read_read_4_stage_61 <= bright_bright_weights_update_0_read_read_4_stage_60;
      bright_bright_weights_update_0_read_read_4_stage_62 <= bright_bright_weights_update_0_read_read_4_stage_61;
      bright_bright_weights_update_0_read_read_4_stage_63 <= bright_bright_weights_update_0_read_read_4_stage_62;
      bright_bright_weights_update_0_read_read_4_stage_64 <= bright_bright_weights_update_0_read_read_4_stage_63;
      bright_bright_weights_update_0_read_read_4_stage_65 <= bright_bright_weights_update_0_read_read_4_stage_64;
      bright_bright_weights_update_0_read_read_4_stage_66 <= bright_bright_weights_update_0_read_read_4_stage_65;
      bright_bright_weights_update_0_read_read_4_stage_67 <= bright_bright_weights_update_0_read_read_4_stage_66;
      bright_bright_weights_update_0_read_read_4_stage_68 <= bright_bright_weights_update_0_read_read_4_stage_67;
      bright_bright_weights_update_0_read_read_4_stage_69 <= bright_bright_weights_update_0_read_read_4_stage_68;
      bright_bright_weights_update_0_read_read_4_stage_70 <= bright_bright_weights_update_0_read_read_4_stage_69;
      bright_bright_weights_update_0_read_read_4_stage_71 <= bright_bright_weights_update_0_read_read_4_stage_70;
      bright_bright_weights_update_0_read_read_4_stage_72 <= bright_bright_weights_update_0_read_read_4_stage_71;
      bright_bright_weights_update_0_read_read_4_stage_73 <= bright_bright_weights_update_0_read_read_4_stage_72;
      bright_bright_weights_update_0_read_read_4_stage_74 <= bright_bright_weights_update_0_read_read_4_stage_73;
      bright_bright_weights_update_0_read_read_4_stage_75 <= bright_bright_weights_update_0_read_read_4_stage_74;
      bright_bright_weights_update_0_read_read_4_stage_76 <= bright_bright_weights_update_0_read_read_4_stage_75;
      bright_bright_weights_update_0_read_read_4_stage_77 <= bright_bright_weights_update_0_read_read_4_stage_76;
      bright_bright_weights_update_0_read_read_4_stage_78 <= bright_bright_weights_update_0_read_read_4_stage_77;
      bright_bright_weights_update_0_read_read_4_stage_79 <= bright_bright_weights_update_0_read_read_4_stage_78;
      bright_bright_weights_update_0_read_read_4_stage_80 <= bright_bright_weights_update_0_read_read_4_stage_79;
      bright_bright_weights_update_0_read_read_4_stage_81 <= bright_bright_weights_update_0_read_read_4_stage_80;
      bright_bright_weights_update_0_read_read_4_stage_82 <= bright_bright_weights_update_0_read_read_4_stage_81;
      bright_bright_weights_update_0_read_read_4_stage_83 <= bright_bright_weights_update_0_read_read_4_stage_82;
      bright_bright_weights_update_0_read_read_4_stage_84 <= bright_bright_weights_update_0_read_read_4_stage_83;
      bright_bright_weights_update_0_read_read_4_stage_85 <= bright_bright_weights_update_0_read_read_4_stage_84;
      bright_bright_weights_update_0_read_read_4_stage_86 <= bright_bright_weights_update_0_read_read_4_stage_85;
      bright_bright_weights_update_0_read_read_4_stage_87 <= bright_bright_weights_update_0_read_read_4_stage_86;
      bright_bright_weights_update_0_read_read_4_stage_88 <= bright_bright_weights_update_0_read_read_4_stage_87;
      bright_bright_weights_update_0_read_read_4_stage_89 <= bright_bright_weights_update_0_read_read_4_stage_88;
      bright_bright_weights_update_0_read_read_4_stage_90 <= bright_bright_weights_update_0_read_read_4_stage_89;
      bright_bright_weights_update_0_read_read_4_stage_91 <= bright_bright_weights_update_0_read_read_4_stage_90;
      bright_bright_weights_update_0_read_read_4_stage_92 <= bright_bright_weights_update_0_read_read_4_stage_91;
      bright_bright_weights_update_0_read_read_4_stage_93 <= bright_bright_weights_update_0_read_read_4_stage_92;
      bright_bright_weights_update_0_read_read_4_stage_94 <= bright_bright_weights_update_0_read_read_4_stage_93;
      bright_bright_weights_update_0_read_read_4_stage_95 <= bright_bright_weights_update_0_read_read_4_stage_94;
      bright_bright_weights_update_0_read_read_4_stage_96 <= bright_bright_weights_update_0_read_read_4_stage_95;
      bright_bright_weights_update_0_read_read_4_stage_97 <= bright_bright_weights_update_0_read_read_4_stage_96;
      bright_bright_weights_update_0_read_read_4_stage_98 <= bright_bright_weights_update_0_read_read_4_stage_97;
      bright_bright_weights_update_0_read_read_4_stage_99 <= bright_bright_weights_update_0_read_read_4_stage_98;
      bright_bright_weights_update_0_read_read_4_stage_100 <= bright_bright_weights_update_0_read_read_4_stage_99;
      bright_bright_weights_update_0_read_read_4_stage_101 <= bright_bright_weights_update_0_read_read_4_stage_100;
      bright_bright_weights_update_0_read_read_4_stage_102 <= bright_bright_weights_update_0_read_read_4_stage_101;
      bright_bright_weights_update_0_read_read_4_stage_103 <= bright_bright_weights_update_0_read_read_4_stage_102;
      bright_bright_weights_update_0_read_read_4_stage_104 <= bright_bright_weights_update_0_read_read_4_stage_103;
      bright_bright_weights_update_0_read_read_4_stage_105 <= bright_bright_weights_update_0_read_read_4_stage_104;
      bright_bright_weights_update_0_read_read_4_stage_106 <= bright_bright_weights_update_0_read_read_4_stage_105;
      bright_bright_weights_update_0_read_read_4_stage_107 <= bright_bright_weights_update_0_read_read_4_stage_106;
      bright_bright_weights_update_0_read_read_4_stage_108 <= bright_bright_weights_update_0_read_read_4_stage_107;
      bright_bright_weights_update_0_read_read_4_stage_109 <= bright_bright_weights_update_0_read_read_4_stage_108;
      bright_bright_weights_update_0_read_read_4_stage_110 <= bright_bright_weights_update_0_read_read_4_stage_109;
      bright_bright_weights_update_0_read_read_4_stage_111 <= bright_bright_weights_update_0_read_read_4_stage_110;
      bright_bright_weights_update_0_read_read_4_stage_112 <= bright_bright_weights_update_0_read_read_4_stage_111;
      bright_bright_weights_update_0_read_read_4_stage_113 <= bright_bright_weights_update_0_read_read_4_stage_112;
      bright_bright_weights_update_0_read_read_4_stage_114 <= bright_bright_weights_update_0_read_read_4_stage_113;
      bright_bright_weights_update_0_read_read_4_stage_115 <= bright_bright_weights_update_0_read_read_4_stage_114;
      bright_bright_weights_update_0_read_read_4_stage_116 <= bright_bright_weights_update_0_read_read_4_stage_115;
      bright_bright_weights_update_0_read_read_4_stage_117 <= bright_bright_weights_update_0_read_read_4_stage_116;
      bright_bright_weights_update_0_read_read_4_stage_118 <= bright_bright_weights_update_0_read_read_4_stage_117;
      bright_bright_weights_update_0_read_read_4_stage_119 <= bright_bright_weights_update_0_read_read_4_stage_118;
      bright_bright_weights_update_0_read_read_4_stage_120 <= bright_bright_weights_update_0_read_read_4_stage_119;
      bright_bright_weights_update_0_read_read_4_stage_121 <= bright_bright_weights_update_0_read_read_4_stage_120;
      bright_bright_weights_update_0_read_read_4_stage_122 <= bright_bright_weights_update_0_read_read_4_stage_121;
      bright_bright_weights_update_0_read_read_4_stage_123 <= bright_bright_weights_update_0_read_read_4_stage_122;
      bright_bright_weights_update_0_read_read_4_stage_124 <= bright_bright_weights_update_0_read_read_4_stage_123;
      bright_bright_weights_update_0_read_read_4_stage_125 <= bright_bright_weights_update_0_read_read_4_stage_124;
      bright_bright_weights_update_0_read_read_4_stage_126 <= bright_bright_weights_update_0_read_read_4_stage_125;
      bright_bright_weights_update_0_read_read_4_stage_127 <= bright_bright_weights_update_0_read_read_4_stage_126;
      bright_bright_weights_update_0_read_read_4_stage_128 <= bright_bright_weights_update_0_read_read_4_stage_127;
      bright_bright_weights_update_0_read_read_4_stage_129 <= bright_bright_weights_update_0_read_read_4_stage_128;
      bright_bright_weights_update_0_read_read_4_stage_130 <= bright_bright_weights_update_0_read_read_4_stage_129;
      bright_bright_weights_update_0_read_read_4_stage_131 <= bright_bright_weights_update_0_read_read_4_stage_130;
      bright_bright_weights_update_0_read_read_4_stage_132 <= bright_bright_weights_update_0_read_read_4_stage_131;
      bright_bright_weights_update_0_read_read_4_stage_133 <= bright_bright_weights_update_0_read_read_4_stage_132;
      bright_bright_weights_update_0_read_read_4_stage_134 <= bright_bright_weights_update_0_read_read_4_stage_133;
      bright_bright_weights_update_0_read_read_4_stage_135 <= bright_bright_weights_update_0_read_read_4_stage_134;
      bright_bright_weights_update_0_read_read_4_stage_136 <= bright_bright_weights_update_0_read_read_4_stage_135;
      bright_bright_weights_update_0_read_read_4_stage_137 <= bright_bright_weights_update_0_read_read_4_stage_136;
      bright_bright_weights_update_0_read_read_4_stage_138 <= bright_bright_weights_update_0_read_read_4_stage_137;
      bright_bright_weights_update_0_read_read_4_stage_139 <= bright_bright_weights_update_0_read_read_4_stage_138;
      bright_bright_weights_update_0_read_read_4_stage_140 <= bright_bright_weights_update_0_read_read_4_stage_139;
      bright_bright_weights_update_0_read_read_4_stage_141 <= bright_bright_weights_update_0_read_read_4_stage_140;
      bright_bright_weights_update_0_read_read_4_stage_142 <= bright_bright_weights_update_0_read_read_4_stage_141;
      bright_bright_weights_update_0_read_read_4_stage_143 <= bright_bright_weights_update_0_read_read_4_stage_142;
      bright_bright_weights_update_0_read_read_4_stage_144 <= bright_bright_weights_update_0_read_read_4_stage_143;
      bright_bright_weights_update_0_read_read_4_stage_145 <= bright_bright_weights_update_0_read_read_4_stage_144;
      bright_bright_weights_update_0_read_read_4_stage_146 <= bright_bright_weights_update_0_read_read_4_stage_145;
      bright_bright_weights_update_0_read_read_4_stage_147 <= bright_bright_weights_update_0_read_read_4_stage_146;
      bright_bright_weights_update_0_read_read_4_stage_148 <= bright_bright_weights_update_0_read_read_4_stage_147;
      bright_bright_weights_update_0_read_read_4_stage_149 <= bright_bright_weights_update_0_read_read_4_stage_148;
      bright_bright_weights_update_0_read_read_4_stage_150 <= bright_bright_weights_update_0_read_read_4_stage_149;
      bright_bright_weights_update_0_read_read_4_stage_151 <= bright_bright_weights_update_0_read_read_4_stage_150;
      bright_bright_weights_update_0_read_read_4_stage_152 <= bright_bright_weights_update_0_read_read_4_stage_151;
      bright_bright_weights_update_0_read_read_4_stage_153 <= bright_bright_weights_update_0_read_read_4_stage_152;
      bright_bright_weights_update_0_read_read_4_stage_154 <= bright_bright_weights_update_0_read_read_4_stage_153;
      bright_bright_weights_update_0_read_read_4_stage_155 <= bright_bright_weights_update_0_read_read_4_stage_154;
      bright_bright_weights_update_0_read_read_4_stage_156 <= bright_bright_weights_update_0_read_read_4_stage_155;
      bright_bright_weights_update_0_read_read_4_stage_157 <= bright_bright_weights_update_0_read_read_4_stage_156;
      bright_bright_weights_update_0_read_read_4_stage_158 <= bright_bright_weights_update_0_read_read_4_stage_157;
      bright_bright_weights_update_0_read_read_4_stage_159 <= bright_bright_weights_update_0_read_read_4_stage_158;
      bright_bright_weights_update_0_read_read_4_stage_160 <= bright_bright_weights_update_0_read_read_4_stage_159;
      bright_bright_weights_update_0_read_read_4_stage_161 <= bright_bright_weights_update_0_read_read_4_stage_160;
      bright_bright_weights_update_0_read_read_4_stage_162 <= bright_bright_weights_update_0_read_read_4_stage_161;
      bright_bright_weights_update_0_read_read_4_stage_163 <= bright_bright_weights_update_0_read_read_4_stage_162;
      bright_bright_weights_update_0_read_read_4_stage_164 <= bright_bright_weights_update_0_read_read_4_stage_163;
      bright_bright_weights_update_0_read_read_4_stage_165 <= bright_bright_weights_update_0_read_read_4_stage_164;
      bright_bright_weights_update_0_read_read_4_stage_166 <= bright_bright_weights_update_0_read_read_4_stage_165;
      bright_bright_weights_update_0_read_read_4_stage_167 <= bright_bright_weights_update_0_read_read_4_stage_166;
      bright_bright_weights_update_0_read_read_4_stage_168 <= bright_bright_weights_update_0_read_read_4_stage_167;
      bright_bright_weights_update_0_read_read_4_stage_169 <= bright_bright_weights_update_0_read_read_4_stage_168;
      bright_bright_weights_update_0_read_read_4_stage_170 <= bright_bright_weights_update_0_read_read_4_stage_169;
      bright_bright_weights_update_0_read_read_4_stage_171 <= bright_bright_weights_update_0_read_read_4_stage_170;
      bright_bright_weights_update_0_read_read_4_stage_172 <= bright_bright_weights_update_0_read_read_4_stage_171;
      bright_bright_weights_update_0_read_read_4_stage_173 <= bright_bright_weights_update_0_read_read_4_stage_172;
      bright_bright_weights_update_0_read_read_4_stage_174 <= bright_bright_weights_update_0_read_read_4_stage_173;
      bright_bright_weights_update_0_read_read_4_stage_175 <= bright_bright_weights_update_0_read_read_4_stage_174;
      bright_bright_weights_update_0_read_read_4_stage_176 <= bright_bright_weights_update_0_read_read_4_stage_175;
      bright_bright_weights_update_0_read_read_4_stage_177 <= bright_bright_weights_update_0_read_read_4_stage_176;
      bright_bright_weights_update_0_read_read_4_stage_178 <= bright_bright_weights_update_0_read_read_4_stage_177;
      bright_bright_weights_update_0_read_read_4_stage_179 <= bright_bright_weights_update_0_read_read_4_stage_178;
      bright_bright_weights_update_0_read_read_4_stage_180 <= bright_bright_weights_update_0_read_read_4_stage_179;
      bright_bright_weights_update_0_read_read_4_stage_181 <= bright_bright_weights_update_0_read_read_4_stage_180;
      bright_weights_update_0_stage_9 <= bright_weights_update_0;
      bright_weights_update_0_stage_10 <= bright_weights_update_0_stage_9;
      bright_weights_update_0_stage_11 <= bright_weights_update_0_stage_10;
      bright_weights_update_0_stage_12 <= bright_weights_update_0_stage_11;
      bright_weights_update_0_stage_13 <= bright_weights_update_0_stage_12;
      bright_weights_update_0_stage_14 <= bright_weights_update_0_stage_13;
      bright_weights_update_0_stage_15 <= bright_weights_update_0_stage_14;
      bright_weights_update_0_stage_16 <= bright_weights_update_0_stage_15;
      bright_weights_update_0_stage_17 <= bright_weights_update_0_stage_16;
      bright_weights_update_0_stage_18 <= bright_weights_update_0_stage_17;
      bright_weights_update_0_stage_19 <= bright_weights_update_0_stage_18;
      bright_weights_update_0_stage_20 <= bright_weights_update_0_stage_19;
      bright_weights_update_0_stage_21 <= bright_weights_update_0_stage_20;
      bright_weights_update_0_stage_22 <= bright_weights_update_0_stage_21;
      bright_weights_update_0_stage_23 <= bright_weights_update_0_stage_22;
      bright_weights_update_0_stage_24 <= bright_weights_update_0_stage_23;
      bright_weights_update_0_stage_25 <= bright_weights_update_0_stage_24;
      bright_weights_update_0_stage_26 <= bright_weights_update_0_stage_25;
      bright_weights_update_0_stage_27 <= bright_weights_update_0_stage_26;
      bright_weights_update_0_stage_28 <= bright_weights_update_0_stage_27;
      bright_weights_update_0_stage_29 <= bright_weights_update_0_stage_28;
      bright_weights_update_0_stage_30 <= bright_weights_update_0_stage_29;
      bright_weights_update_0_stage_31 <= bright_weights_update_0_stage_30;
      bright_weights_update_0_stage_32 <= bright_weights_update_0_stage_31;
      bright_weights_update_0_stage_33 <= bright_weights_update_0_stage_32;
      bright_weights_update_0_stage_34 <= bright_weights_update_0_stage_33;
      bright_weights_update_0_stage_35 <= bright_weights_update_0_stage_34;
      bright_weights_update_0_stage_36 <= bright_weights_update_0_stage_35;
      bright_weights_update_0_stage_37 <= bright_weights_update_0_stage_36;
      bright_weights_update_0_stage_38 <= bright_weights_update_0_stage_37;
      bright_weights_update_0_stage_39 <= bright_weights_update_0_stage_38;
      bright_weights_update_0_stage_40 <= bright_weights_update_0_stage_39;
      bright_weights_update_0_stage_41 <= bright_weights_update_0_stage_40;
      bright_weights_update_0_stage_42 <= bright_weights_update_0_stage_41;
      bright_weights_update_0_stage_43 <= bright_weights_update_0_stage_42;
      bright_weights_update_0_stage_44 <= bright_weights_update_0_stage_43;
      bright_weights_update_0_stage_45 <= bright_weights_update_0_stage_44;
      bright_weights_update_0_stage_46 <= bright_weights_update_0_stage_45;
      bright_weights_update_0_stage_47 <= bright_weights_update_0_stage_46;
      bright_weights_update_0_stage_48 <= bright_weights_update_0_stage_47;
      bright_weights_update_0_stage_49 <= bright_weights_update_0_stage_48;
      bright_weights_update_0_stage_50 <= bright_weights_update_0_stage_49;
      bright_weights_update_0_stage_51 <= bright_weights_update_0_stage_50;
      bright_weights_update_0_stage_52 <= bright_weights_update_0_stage_51;
      bright_weights_update_0_stage_53 <= bright_weights_update_0_stage_52;
      bright_weights_update_0_stage_54 <= bright_weights_update_0_stage_53;
      bright_weights_update_0_stage_55 <= bright_weights_update_0_stage_54;
      bright_weights_update_0_stage_56 <= bright_weights_update_0_stage_55;
      bright_weights_update_0_stage_57 <= bright_weights_update_0_stage_56;
      bright_weights_update_0_stage_58 <= bright_weights_update_0_stage_57;
      bright_weights_update_0_stage_59 <= bright_weights_update_0_stage_58;
      bright_weights_update_0_stage_60 <= bright_weights_update_0_stage_59;
      bright_weights_update_0_stage_61 <= bright_weights_update_0_stage_60;
      bright_weights_update_0_stage_62 <= bright_weights_update_0_stage_61;
      bright_weights_update_0_stage_63 <= bright_weights_update_0_stage_62;
      bright_weights_update_0_stage_64 <= bright_weights_update_0_stage_63;
      bright_weights_update_0_stage_65 <= bright_weights_update_0_stage_64;
      bright_weights_update_0_stage_66 <= bright_weights_update_0_stage_65;
      bright_weights_update_0_stage_67 <= bright_weights_update_0_stage_66;
      bright_weights_update_0_stage_68 <= bright_weights_update_0_stage_67;
      bright_weights_update_0_stage_69 <= bright_weights_update_0_stage_68;
      bright_weights_update_0_stage_70 <= bright_weights_update_0_stage_69;
      bright_weights_update_0_stage_71 <= bright_weights_update_0_stage_70;
      bright_weights_update_0_stage_72 <= bright_weights_update_0_stage_71;
      bright_weights_update_0_stage_73 <= bright_weights_update_0_stage_72;
      bright_weights_update_0_stage_74 <= bright_weights_update_0_stage_73;
      bright_weights_update_0_stage_75 <= bright_weights_update_0_stage_74;
      bright_weights_update_0_stage_76 <= bright_weights_update_0_stage_75;
      bright_weights_update_0_stage_77 <= bright_weights_update_0_stage_76;
      bright_weights_update_0_stage_78 <= bright_weights_update_0_stage_77;
      bright_weights_update_0_stage_79 <= bright_weights_update_0_stage_78;
      bright_weights_update_0_stage_80 <= bright_weights_update_0_stage_79;
      bright_weights_update_0_stage_81 <= bright_weights_update_0_stage_80;
      bright_weights_update_0_stage_82 <= bright_weights_update_0_stage_81;
      bright_weights_update_0_stage_83 <= bright_weights_update_0_stage_82;
      bright_weights_update_0_stage_84 <= bright_weights_update_0_stage_83;
      bright_weights_update_0_stage_85 <= bright_weights_update_0_stage_84;
      bright_weights_update_0_stage_86 <= bright_weights_update_0_stage_85;
      bright_weights_update_0_stage_87 <= bright_weights_update_0_stage_86;
      bright_weights_update_0_stage_88 <= bright_weights_update_0_stage_87;
      bright_weights_update_0_stage_89 <= bright_weights_update_0_stage_88;
      bright_weights_update_0_stage_90 <= bright_weights_update_0_stage_89;
      bright_weights_update_0_stage_91 <= bright_weights_update_0_stage_90;
      bright_weights_update_0_stage_92 <= bright_weights_update_0_stage_91;
      bright_weights_update_0_stage_93 <= bright_weights_update_0_stage_92;
      bright_weights_update_0_stage_94 <= bright_weights_update_0_stage_93;
      bright_weights_update_0_stage_95 <= bright_weights_update_0_stage_94;
      bright_weights_update_0_stage_96 <= bright_weights_update_0_stage_95;
      bright_weights_update_0_stage_97 <= bright_weights_update_0_stage_96;
      bright_weights_update_0_stage_98 <= bright_weights_update_0_stage_97;
      bright_weights_update_0_stage_99 <= bright_weights_update_0_stage_98;
      bright_weights_update_0_stage_100 <= bright_weights_update_0_stage_99;
      bright_weights_update_0_stage_101 <= bright_weights_update_0_stage_100;
      bright_weights_update_0_stage_102 <= bright_weights_update_0_stage_101;
      bright_weights_update_0_stage_103 <= bright_weights_update_0_stage_102;
      bright_weights_update_0_stage_104 <= bright_weights_update_0_stage_103;
      bright_weights_update_0_stage_105 <= bright_weights_update_0_stage_104;
      bright_weights_update_0_stage_106 <= bright_weights_update_0_stage_105;
      bright_weights_update_0_stage_107 <= bright_weights_update_0_stage_106;
      bright_weights_update_0_stage_108 <= bright_weights_update_0_stage_107;
      bright_weights_update_0_stage_109 <= bright_weights_update_0_stage_108;
      bright_weights_update_0_stage_110 <= bright_weights_update_0_stage_109;
      bright_weights_update_0_stage_111 <= bright_weights_update_0_stage_110;
      bright_weights_update_0_stage_112 <= bright_weights_update_0_stage_111;
      bright_weights_update_0_stage_113 <= bright_weights_update_0_stage_112;
      bright_weights_update_0_stage_114 <= bright_weights_update_0_stage_113;
      bright_weights_update_0_stage_115 <= bright_weights_update_0_stage_114;
      bright_weights_update_0_stage_116 <= bright_weights_update_0_stage_115;
      bright_weights_update_0_stage_117 <= bright_weights_update_0_stage_116;
      bright_weights_update_0_stage_118 <= bright_weights_update_0_stage_117;
      bright_weights_update_0_stage_119 <= bright_weights_update_0_stage_118;
      bright_weights_update_0_stage_120 <= bright_weights_update_0_stage_119;
      bright_weights_update_0_stage_121 <= bright_weights_update_0_stage_120;
      bright_weights_update_0_stage_122 <= bright_weights_update_0_stage_121;
      bright_weights_update_0_stage_123 <= bright_weights_update_0_stage_122;
      bright_weights_update_0_stage_124 <= bright_weights_update_0_stage_123;
      bright_weights_update_0_stage_125 <= bright_weights_update_0_stage_124;
      bright_weights_update_0_stage_126 <= bright_weights_update_0_stage_125;
      bright_weights_update_0_stage_127 <= bright_weights_update_0_stage_126;
      bright_weights_update_0_stage_128 <= bright_weights_update_0_stage_127;
      bright_weights_update_0_stage_129 <= bright_weights_update_0_stage_128;
      bright_weights_update_0_stage_130 <= bright_weights_update_0_stage_129;
      bright_weights_update_0_stage_131 <= bright_weights_update_0_stage_130;
      bright_weights_update_0_stage_132 <= bright_weights_update_0_stage_131;
      bright_weights_update_0_stage_133 <= bright_weights_update_0_stage_132;
      bright_weights_update_0_stage_134 <= bright_weights_update_0_stage_133;
      bright_weights_update_0_stage_135 <= bright_weights_update_0_stage_134;
      bright_weights_update_0_stage_136 <= bright_weights_update_0_stage_135;
      bright_weights_update_0_stage_137 <= bright_weights_update_0_stage_136;
      bright_weights_update_0_stage_138 <= bright_weights_update_0_stage_137;
      bright_weights_update_0_stage_139 <= bright_weights_update_0_stage_138;
      bright_weights_update_0_stage_140 <= bright_weights_update_0_stage_139;
      bright_weights_update_0_stage_141 <= bright_weights_update_0_stage_140;
      bright_weights_update_0_stage_142 <= bright_weights_update_0_stage_141;
      bright_weights_update_0_stage_143 <= bright_weights_update_0_stage_142;
      bright_weights_update_0_stage_144 <= bright_weights_update_0_stage_143;
      bright_weights_update_0_stage_145 <= bright_weights_update_0_stage_144;
      bright_weights_update_0_stage_146 <= bright_weights_update_0_stage_145;
      bright_weights_update_0_stage_147 <= bright_weights_update_0_stage_146;
      bright_weights_update_0_stage_148 <= bright_weights_update_0_stage_147;
      bright_weights_update_0_stage_149 <= bright_weights_update_0_stage_148;
      bright_weights_update_0_stage_150 <= bright_weights_update_0_stage_149;
      bright_weights_update_0_stage_151 <= bright_weights_update_0_stage_150;
      bright_weights_update_0_stage_152 <= bright_weights_update_0_stage_151;
      bright_weights_update_0_stage_153 <= bright_weights_update_0_stage_152;
      bright_weights_update_0_stage_154 <= bright_weights_update_0_stage_153;
      bright_weights_update_0_stage_155 <= bright_weights_update_0_stage_154;
      bright_weights_update_0_stage_156 <= bright_weights_update_0_stage_155;
      bright_weights_update_0_stage_157 <= bright_weights_update_0_stage_156;
      bright_weights_update_0_stage_158 <= bright_weights_update_0_stage_157;
      bright_weights_update_0_stage_159 <= bright_weights_update_0_stage_158;
      bright_weights_update_0_stage_160 <= bright_weights_update_0_stage_159;
      bright_weights_update_0_stage_161 <= bright_weights_update_0_stage_160;
      bright_weights_update_0_stage_162 <= bright_weights_update_0_stage_161;
      bright_weights_update_0_stage_163 <= bright_weights_update_0_stage_162;
      bright_weights_update_0_stage_164 <= bright_weights_update_0_stage_163;
      bright_weights_update_0_stage_165 <= bright_weights_update_0_stage_164;
      bright_weights_update_0_stage_166 <= bright_weights_update_0_stage_165;
      bright_weights_update_0_stage_167 <= bright_weights_update_0_stage_166;
      bright_weights_update_0_stage_168 <= bright_weights_update_0_stage_167;
      bright_weights_update_0_stage_169 <= bright_weights_update_0_stage_168;
      bright_weights_update_0_stage_170 <= bright_weights_update_0_stage_169;
      bright_weights_update_0_stage_171 <= bright_weights_update_0_stage_170;
      bright_weights_update_0_stage_172 <= bright_weights_update_0_stage_171;
      bright_weights_update_0_stage_173 <= bright_weights_update_0_stage_172;
      bright_weights_update_0_stage_174 <= bright_weights_update_0_stage_173;
      bright_weights_update_0_stage_175 <= bright_weights_update_0_stage_174;
      bright_weights_update_0_stage_176 <= bright_weights_update_0_stage_175;
      bright_weights_update_0_stage_177 <= bright_weights_update_0_stage_176;
      bright_weights_update_0_stage_178 <= bright_weights_update_0_stage_177;
      bright_weights_update_0_stage_179 <= bright_weights_update_0_stage_178;
      bright_weights_update_0_stage_180 <= bright_weights_update_0_stage_179;
      bright_weights_update_0_stage_181 <= bright_weights_update_0_stage_180;
      bright_weights_bright_weights_update_0_write_write_5_stage_10 <= bright_weights_bright_weights_update_0_write_write_5;
      bright_weights_bright_weights_update_0_write_write_5_stage_11 <= bright_weights_bright_weights_update_0_write_write_5_stage_10;
      bright_weights_bright_weights_update_0_write_write_5_stage_12 <= bright_weights_bright_weights_update_0_write_write_5_stage_11;
      bright_weights_bright_weights_update_0_write_write_5_stage_13 <= bright_weights_bright_weights_update_0_write_write_5_stage_12;
      bright_weights_bright_weights_update_0_write_write_5_stage_14 <= bright_weights_bright_weights_update_0_write_write_5_stage_13;
      bright_weights_bright_weights_update_0_write_write_5_stage_15 <= bright_weights_bright_weights_update_0_write_write_5_stage_14;
      bright_weights_bright_weights_update_0_write_write_5_stage_16 <= bright_weights_bright_weights_update_0_write_write_5_stage_15;
      bright_weights_bright_weights_update_0_write_write_5_stage_17 <= bright_weights_bright_weights_update_0_write_write_5_stage_16;
      bright_weights_bright_weights_update_0_write_write_5_stage_18 <= bright_weights_bright_weights_update_0_write_write_5_stage_17;
      bright_weights_bright_weights_update_0_write_write_5_stage_19 <= bright_weights_bright_weights_update_0_write_write_5_stage_18;
      bright_weights_bright_weights_update_0_write_write_5_stage_20 <= bright_weights_bright_weights_update_0_write_write_5_stage_19;
      bright_weights_bright_weights_update_0_write_write_5_stage_21 <= bright_weights_bright_weights_update_0_write_write_5_stage_20;
      bright_weights_bright_weights_update_0_write_write_5_stage_22 <= bright_weights_bright_weights_update_0_write_write_5_stage_21;
      bright_weights_bright_weights_update_0_write_write_5_stage_23 <= bright_weights_bright_weights_update_0_write_write_5_stage_22;
      bright_weights_bright_weights_update_0_write_write_5_stage_24 <= bright_weights_bright_weights_update_0_write_write_5_stage_23;
      bright_weights_bright_weights_update_0_write_write_5_stage_25 <= bright_weights_bright_weights_update_0_write_write_5_stage_24;
      bright_weights_bright_weights_update_0_write_write_5_stage_26 <= bright_weights_bright_weights_update_0_write_write_5_stage_25;
      bright_weights_bright_weights_update_0_write_write_5_stage_27 <= bright_weights_bright_weights_update_0_write_write_5_stage_26;
      bright_weights_bright_weights_update_0_write_write_5_stage_28 <= bright_weights_bright_weights_update_0_write_write_5_stage_27;
      bright_weights_bright_weights_update_0_write_write_5_stage_29 <= bright_weights_bright_weights_update_0_write_write_5_stage_28;
      bright_weights_bright_weights_update_0_write_write_5_stage_30 <= bright_weights_bright_weights_update_0_write_write_5_stage_29;
      bright_weights_bright_weights_update_0_write_write_5_stage_31 <= bright_weights_bright_weights_update_0_write_write_5_stage_30;
      bright_weights_bright_weights_update_0_write_write_5_stage_32 <= bright_weights_bright_weights_update_0_write_write_5_stage_31;
      bright_weights_bright_weights_update_0_write_write_5_stage_33 <= bright_weights_bright_weights_update_0_write_write_5_stage_32;
      bright_weights_bright_weights_update_0_write_write_5_stage_34 <= bright_weights_bright_weights_update_0_write_write_5_stage_33;
      bright_weights_bright_weights_update_0_write_write_5_stage_35 <= bright_weights_bright_weights_update_0_write_write_5_stage_34;
      bright_weights_bright_weights_update_0_write_write_5_stage_36 <= bright_weights_bright_weights_update_0_write_write_5_stage_35;
      bright_weights_bright_weights_update_0_write_write_5_stage_37 <= bright_weights_bright_weights_update_0_write_write_5_stage_36;
      bright_weights_bright_weights_update_0_write_write_5_stage_38 <= bright_weights_bright_weights_update_0_write_write_5_stage_37;
      bright_weights_bright_weights_update_0_write_write_5_stage_39 <= bright_weights_bright_weights_update_0_write_write_5_stage_38;
      bright_weights_bright_weights_update_0_write_write_5_stage_40 <= bright_weights_bright_weights_update_0_write_write_5_stage_39;
      bright_weights_bright_weights_update_0_write_write_5_stage_41 <= bright_weights_bright_weights_update_0_write_write_5_stage_40;
      bright_weights_bright_weights_update_0_write_write_5_stage_42 <= bright_weights_bright_weights_update_0_write_write_5_stage_41;
      bright_weights_bright_weights_update_0_write_write_5_stage_43 <= bright_weights_bright_weights_update_0_write_write_5_stage_42;
      bright_weights_bright_weights_update_0_write_write_5_stage_44 <= bright_weights_bright_weights_update_0_write_write_5_stage_43;
      bright_weights_bright_weights_update_0_write_write_5_stage_45 <= bright_weights_bright_weights_update_0_write_write_5_stage_44;
      bright_weights_bright_weights_update_0_write_write_5_stage_46 <= bright_weights_bright_weights_update_0_write_write_5_stage_45;
      bright_weights_bright_weights_update_0_write_write_5_stage_47 <= bright_weights_bright_weights_update_0_write_write_5_stage_46;
      bright_weights_bright_weights_update_0_write_write_5_stage_48 <= bright_weights_bright_weights_update_0_write_write_5_stage_47;
      bright_weights_bright_weights_update_0_write_write_5_stage_49 <= bright_weights_bright_weights_update_0_write_write_5_stage_48;
      bright_weights_bright_weights_update_0_write_write_5_stage_50 <= bright_weights_bright_weights_update_0_write_write_5_stage_49;
      bright_weights_bright_weights_update_0_write_write_5_stage_51 <= bright_weights_bright_weights_update_0_write_write_5_stage_50;
      bright_weights_bright_weights_update_0_write_write_5_stage_52 <= bright_weights_bright_weights_update_0_write_write_5_stage_51;
      bright_weights_bright_weights_update_0_write_write_5_stage_53 <= bright_weights_bright_weights_update_0_write_write_5_stage_52;
      bright_weights_bright_weights_update_0_write_write_5_stage_54 <= bright_weights_bright_weights_update_0_write_write_5_stage_53;
      bright_weights_bright_weights_update_0_write_write_5_stage_55 <= bright_weights_bright_weights_update_0_write_write_5_stage_54;
      bright_weights_bright_weights_update_0_write_write_5_stage_56 <= bright_weights_bright_weights_update_0_write_write_5_stage_55;
      bright_weights_bright_weights_update_0_write_write_5_stage_57 <= bright_weights_bright_weights_update_0_write_write_5_stage_56;
      bright_weights_bright_weights_update_0_write_write_5_stage_58 <= bright_weights_bright_weights_update_0_write_write_5_stage_57;
      bright_weights_bright_weights_update_0_write_write_5_stage_59 <= bright_weights_bright_weights_update_0_write_write_5_stage_58;
      bright_weights_bright_weights_update_0_write_write_5_stage_60 <= bright_weights_bright_weights_update_0_write_write_5_stage_59;
      bright_weights_bright_weights_update_0_write_write_5_stage_61 <= bright_weights_bright_weights_update_0_write_write_5_stage_60;
      bright_weights_bright_weights_update_0_write_write_5_stage_62 <= bright_weights_bright_weights_update_0_write_write_5_stage_61;
      bright_weights_bright_weights_update_0_write_write_5_stage_63 <= bright_weights_bright_weights_update_0_write_write_5_stage_62;
      bright_weights_bright_weights_update_0_write_write_5_stage_64 <= bright_weights_bright_weights_update_0_write_write_5_stage_63;
      bright_weights_bright_weights_update_0_write_write_5_stage_65 <= bright_weights_bright_weights_update_0_write_write_5_stage_64;
      bright_weights_bright_weights_update_0_write_write_5_stage_66 <= bright_weights_bright_weights_update_0_write_write_5_stage_65;
      bright_weights_bright_weights_update_0_write_write_5_stage_67 <= bright_weights_bright_weights_update_0_write_write_5_stage_66;
      bright_weights_bright_weights_update_0_write_write_5_stage_68 <= bright_weights_bright_weights_update_0_write_write_5_stage_67;
      bright_weights_bright_weights_update_0_write_write_5_stage_69 <= bright_weights_bright_weights_update_0_write_write_5_stage_68;
      bright_weights_bright_weights_update_0_write_write_5_stage_70 <= bright_weights_bright_weights_update_0_write_write_5_stage_69;
      bright_weights_bright_weights_update_0_write_write_5_stage_71 <= bright_weights_bright_weights_update_0_write_write_5_stage_70;
      bright_weights_bright_weights_update_0_write_write_5_stage_72 <= bright_weights_bright_weights_update_0_write_write_5_stage_71;
      bright_weights_bright_weights_update_0_write_write_5_stage_73 <= bright_weights_bright_weights_update_0_write_write_5_stage_72;
      bright_weights_bright_weights_update_0_write_write_5_stage_74 <= bright_weights_bright_weights_update_0_write_write_5_stage_73;
      bright_weights_bright_weights_update_0_write_write_5_stage_75 <= bright_weights_bright_weights_update_0_write_write_5_stage_74;
      bright_weights_bright_weights_update_0_write_write_5_stage_76 <= bright_weights_bright_weights_update_0_write_write_5_stage_75;
      bright_weights_bright_weights_update_0_write_write_5_stage_77 <= bright_weights_bright_weights_update_0_write_write_5_stage_76;
      bright_weights_bright_weights_update_0_write_write_5_stage_78 <= bright_weights_bright_weights_update_0_write_write_5_stage_77;
      bright_weights_bright_weights_update_0_write_write_5_stage_79 <= bright_weights_bright_weights_update_0_write_write_5_stage_78;
      bright_weights_bright_weights_update_0_write_write_5_stage_80 <= bright_weights_bright_weights_update_0_write_write_5_stage_79;
      bright_weights_bright_weights_update_0_write_write_5_stage_81 <= bright_weights_bright_weights_update_0_write_write_5_stage_80;
      bright_weights_bright_weights_update_0_write_write_5_stage_82 <= bright_weights_bright_weights_update_0_write_write_5_stage_81;
      bright_weights_bright_weights_update_0_write_write_5_stage_83 <= bright_weights_bright_weights_update_0_write_write_5_stage_82;
      bright_weights_bright_weights_update_0_write_write_5_stage_84 <= bright_weights_bright_weights_update_0_write_write_5_stage_83;
      bright_weights_bright_weights_update_0_write_write_5_stage_85 <= bright_weights_bright_weights_update_0_write_write_5_stage_84;
      bright_weights_bright_weights_update_0_write_write_5_stage_86 <= bright_weights_bright_weights_update_0_write_write_5_stage_85;
      bright_weights_bright_weights_update_0_write_write_5_stage_87 <= bright_weights_bright_weights_update_0_write_write_5_stage_86;
      bright_weights_bright_weights_update_0_write_write_5_stage_88 <= bright_weights_bright_weights_update_0_write_write_5_stage_87;
      bright_weights_bright_weights_update_0_write_write_5_stage_89 <= bright_weights_bright_weights_update_0_write_write_5_stage_88;
      bright_weights_bright_weights_update_0_write_write_5_stage_90 <= bright_weights_bright_weights_update_0_write_write_5_stage_89;
      bright_weights_bright_weights_update_0_write_write_5_stage_91 <= bright_weights_bright_weights_update_0_write_write_5_stage_90;
      bright_weights_bright_weights_update_0_write_write_5_stage_92 <= bright_weights_bright_weights_update_0_write_write_5_stage_91;
      bright_weights_bright_weights_update_0_write_write_5_stage_93 <= bright_weights_bright_weights_update_0_write_write_5_stage_92;
      bright_weights_bright_weights_update_0_write_write_5_stage_94 <= bright_weights_bright_weights_update_0_write_write_5_stage_93;
      bright_weights_bright_weights_update_0_write_write_5_stage_95 <= bright_weights_bright_weights_update_0_write_write_5_stage_94;
      bright_weights_bright_weights_update_0_write_write_5_stage_96 <= bright_weights_bright_weights_update_0_write_write_5_stage_95;
      bright_weights_bright_weights_update_0_write_write_5_stage_97 <= bright_weights_bright_weights_update_0_write_write_5_stage_96;
      bright_weights_bright_weights_update_0_write_write_5_stage_98 <= bright_weights_bright_weights_update_0_write_write_5_stage_97;
      bright_weights_bright_weights_update_0_write_write_5_stage_99 <= bright_weights_bright_weights_update_0_write_write_5_stage_98;
      bright_weights_bright_weights_update_0_write_write_5_stage_100 <= bright_weights_bright_weights_update_0_write_write_5_stage_99;
      bright_weights_bright_weights_update_0_write_write_5_stage_101 <= bright_weights_bright_weights_update_0_write_write_5_stage_100;
      bright_weights_bright_weights_update_0_write_write_5_stage_102 <= bright_weights_bright_weights_update_0_write_write_5_stage_101;
      bright_weights_bright_weights_update_0_write_write_5_stage_103 <= bright_weights_bright_weights_update_0_write_write_5_stage_102;
      bright_weights_bright_weights_update_0_write_write_5_stage_104 <= bright_weights_bright_weights_update_0_write_write_5_stage_103;
      bright_weights_bright_weights_update_0_write_write_5_stage_105 <= bright_weights_bright_weights_update_0_write_write_5_stage_104;
      bright_weights_bright_weights_update_0_write_write_5_stage_106 <= bright_weights_bright_weights_update_0_write_write_5_stage_105;
      bright_weights_bright_weights_update_0_write_write_5_stage_107 <= bright_weights_bright_weights_update_0_write_write_5_stage_106;
      bright_weights_bright_weights_update_0_write_write_5_stage_108 <= bright_weights_bright_weights_update_0_write_write_5_stage_107;
      bright_weights_bright_weights_update_0_write_write_5_stage_109 <= bright_weights_bright_weights_update_0_write_write_5_stage_108;
      bright_weights_bright_weights_update_0_write_write_5_stage_110 <= bright_weights_bright_weights_update_0_write_write_5_stage_109;
      bright_weights_bright_weights_update_0_write_write_5_stage_111 <= bright_weights_bright_weights_update_0_write_write_5_stage_110;
      bright_weights_bright_weights_update_0_write_write_5_stage_112 <= bright_weights_bright_weights_update_0_write_write_5_stage_111;
      bright_weights_bright_weights_update_0_write_write_5_stage_113 <= bright_weights_bright_weights_update_0_write_write_5_stage_112;
      bright_weights_bright_weights_update_0_write_write_5_stage_114 <= bright_weights_bright_weights_update_0_write_write_5_stage_113;
      bright_weights_bright_weights_update_0_write_write_5_stage_115 <= bright_weights_bright_weights_update_0_write_write_5_stage_114;
      bright_weights_bright_weights_update_0_write_write_5_stage_116 <= bright_weights_bright_weights_update_0_write_write_5_stage_115;
      bright_weights_bright_weights_update_0_write_write_5_stage_117 <= bright_weights_bright_weights_update_0_write_write_5_stage_116;
      bright_weights_bright_weights_update_0_write_write_5_stage_118 <= bright_weights_bright_weights_update_0_write_write_5_stage_117;
      bright_weights_bright_weights_update_0_write_write_5_stage_119 <= bright_weights_bright_weights_update_0_write_write_5_stage_118;
      bright_weights_bright_weights_update_0_write_write_5_stage_120 <= bright_weights_bright_weights_update_0_write_write_5_stage_119;
      bright_weights_bright_weights_update_0_write_write_5_stage_121 <= bright_weights_bright_weights_update_0_write_write_5_stage_120;
      bright_weights_bright_weights_update_0_write_write_5_stage_122 <= bright_weights_bright_weights_update_0_write_write_5_stage_121;
      bright_weights_bright_weights_update_0_write_write_5_stage_123 <= bright_weights_bright_weights_update_0_write_write_5_stage_122;
      bright_weights_bright_weights_update_0_write_write_5_stage_124 <= bright_weights_bright_weights_update_0_write_write_5_stage_123;
      bright_weights_bright_weights_update_0_write_write_5_stage_125 <= bright_weights_bright_weights_update_0_write_write_5_stage_124;
      bright_weights_bright_weights_update_0_write_write_5_stage_126 <= bright_weights_bright_weights_update_0_write_write_5_stage_125;
      bright_weights_bright_weights_update_0_write_write_5_stage_127 <= bright_weights_bright_weights_update_0_write_write_5_stage_126;
      bright_weights_bright_weights_update_0_write_write_5_stage_128 <= bright_weights_bright_weights_update_0_write_write_5_stage_127;
      bright_weights_bright_weights_update_0_write_write_5_stage_129 <= bright_weights_bright_weights_update_0_write_write_5_stage_128;
      bright_weights_bright_weights_update_0_write_write_5_stage_130 <= bright_weights_bright_weights_update_0_write_write_5_stage_129;
      bright_weights_bright_weights_update_0_write_write_5_stage_131 <= bright_weights_bright_weights_update_0_write_write_5_stage_130;
      bright_weights_bright_weights_update_0_write_write_5_stage_132 <= bright_weights_bright_weights_update_0_write_write_5_stage_131;
      bright_weights_bright_weights_update_0_write_write_5_stage_133 <= bright_weights_bright_weights_update_0_write_write_5_stage_132;
      bright_weights_bright_weights_update_0_write_write_5_stage_134 <= bright_weights_bright_weights_update_0_write_write_5_stage_133;
      bright_weights_bright_weights_update_0_write_write_5_stage_135 <= bright_weights_bright_weights_update_0_write_write_5_stage_134;
      bright_weights_bright_weights_update_0_write_write_5_stage_136 <= bright_weights_bright_weights_update_0_write_write_5_stage_135;
      bright_weights_bright_weights_update_0_write_write_5_stage_137 <= bright_weights_bright_weights_update_0_write_write_5_stage_136;
      bright_weights_bright_weights_update_0_write_write_5_stage_138 <= bright_weights_bright_weights_update_0_write_write_5_stage_137;
      bright_weights_bright_weights_update_0_write_write_5_stage_139 <= bright_weights_bright_weights_update_0_write_write_5_stage_138;
      bright_weights_bright_weights_update_0_write_write_5_stage_140 <= bright_weights_bright_weights_update_0_write_write_5_stage_139;
      bright_weights_bright_weights_update_0_write_write_5_stage_141 <= bright_weights_bright_weights_update_0_write_write_5_stage_140;
      bright_weights_bright_weights_update_0_write_write_5_stage_142 <= bright_weights_bright_weights_update_0_write_write_5_stage_141;
      bright_weights_bright_weights_update_0_write_write_5_stage_143 <= bright_weights_bright_weights_update_0_write_write_5_stage_142;
      bright_weights_bright_weights_update_0_write_write_5_stage_144 <= bright_weights_bright_weights_update_0_write_write_5_stage_143;
      bright_weights_bright_weights_update_0_write_write_5_stage_145 <= bright_weights_bright_weights_update_0_write_write_5_stage_144;
      bright_weights_bright_weights_update_0_write_write_5_stage_146 <= bright_weights_bright_weights_update_0_write_write_5_stage_145;
      bright_weights_bright_weights_update_0_write_write_5_stage_147 <= bright_weights_bright_weights_update_0_write_write_5_stage_146;
      bright_weights_bright_weights_update_0_write_write_5_stage_148 <= bright_weights_bright_weights_update_0_write_write_5_stage_147;
      bright_weights_bright_weights_update_0_write_write_5_stage_149 <= bright_weights_bright_weights_update_0_write_write_5_stage_148;
      bright_weights_bright_weights_update_0_write_write_5_stage_150 <= bright_weights_bright_weights_update_0_write_write_5_stage_149;
      bright_weights_bright_weights_update_0_write_write_5_stage_151 <= bright_weights_bright_weights_update_0_write_write_5_stage_150;
      bright_weights_bright_weights_update_0_write_write_5_stage_152 <= bright_weights_bright_weights_update_0_write_write_5_stage_151;
      bright_weights_bright_weights_update_0_write_write_5_stage_153 <= bright_weights_bright_weights_update_0_write_write_5_stage_152;
      bright_weights_bright_weights_update_0_write_write_5_stage_154 <= bright_weights_bright_weights_update_0_write_write_5_stage_153;
      bright_weights_bright_weights_update_0_write_write_5_stage_155 <= bright_weights_bright_weights_update_0_write_write_5_stage_154;
      bright_weights_bright_weights_update_0_write_write_5_stage_156 <= bright_weights_bright_weights_update_0_write_write_5_stage_155;
      bright_weights_bright_weights_update_0_write_write_5_stage_157 <= bright_weights_bright_weights_update_0_write_write_5_stage_156;
      bright_weights_bright_weights_update_0_write_write_5_stage_158 <= bright_weights_bright_weights_update_0_write_write_5_stage_157;
      bright_weights_bright_weights_update_0_write_write_5_stage_159 <= bright_weights_bright_weights_update_0_write_write_5_stage_158;
      bright_weights_bright_weights_update_0_write_write_5_stage_160 <= bright_weights_bright_weights_update_0_write_write_5_stage_159;
      bright_weights_bright_weights_update_0_write_write_5_stage_161 <= bright_weights_bright_weights_update_0_write_write_5_stage_160;
      bright_weights_bright_weights_update_0_write_write_5_stage_162 <= bright_weights_bright_weights_update_0_write_write_5_stage_161;
      bright_weights_bright_weights_update_0_write_write_5_stage_163 <= bright_weights_bright_weights_update_0_write_write_5_stage_162;
      bright_weights_bright_weights_update_0_write_write_5_stage_164 <= bright_weights_bright_weights_update_0_write_write_5_stage_163;
      bright_weights_bright_weights_update_0_write_write_5_stage_165 <= bright_weights_bright_weights_update_0_write_write_5_stage_164;
      bright_weights_bright_weights_update_0_write_write_5_stage_166 <= bright_weights_bright_weights_update_0_write_write_5_stage_165;
      bright_weights_bright_weights_update_0_write_write_5_stage_167 <= bright_weights_bright_weights_update_0_write_write_5_stage_166;
      bright_weights_bright_weights_update_0_write_write_5_stage_168 <= bright_weights_bright_weights_update_0_write_write_5_stage_167;
      bright_weights_bright_weights_update_0_write_write_5_stage_169 <= bright_weights_bright_weights_update_0_write_write_5_stage_168;
      bright_weights_bright_weights_update_0_write_write_5_stage_170 <= bright_weights_bright_weights_update_0_write_write_5_stage_169;
      bright_weights_bright_weights_update_0_write_write_5_stage_171 <= bright_weights_bright_weights_update_0_write_write_5_stage_170;
      bright_weights_bright_weights_update_0_write_write_5_stage_172 <= bright_weights_bright_weights_update_0_write_write_5_stage_171;
      bright_weights_bright_weights_update_0_write_write_5_stage_173 <= bright_weights_bright_weights_update_0_write_write_5_stage_172;
      bright_weights_bright_weights_update_0_write_write_5_stage_174 <= bright_weights_bright_weights_update_0_write_write_5_stage_173;
      bright_weights_bright_weights_update_0_write_write_5_stage_175 <= bright_weights_bright_weights_update_0_write_write_5_stage_174;
      bright_weights_bright_weights_update_0_write_write_5_stage_176 <= bright_weights_bright_weights_update_0_write_write_5_stage_175;
      bright_weights_bright_weights_update_0_write_write_5_stage_177 <= bright_weights_bright_weights_update_0_write_write_5_stage_176;
      bright_weights_bright_weights_update_0_write_write_5_stage_178 <= bright_weights_bright_weights_update_0_write_write_5_stage_177;
      bright_weights_bright_weights_update_0_write_write_5_stage_179 <= bright_weights_bright_weights_update_0_write_write_5_stage_178;
      bright_weights_bright_weights_update_0_write_write_5_stage_180 <= bright_weights_bright_weights_update_0_write_write_5_stage_179;
      bright_weights_bright_weights_update_0_write_write_5_stage_181 <= bright_weights_bright_weights_update_0_write_write_5_stage_180;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_85 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_86 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_85;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_87 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_86;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_88 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_87;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_89 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_88;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_90 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_89;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_91 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_90;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_92 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_91;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_93 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_92;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_94 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_93;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_95 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_94;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_96 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_95;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_97 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_96;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_98 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_97;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_99 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_98;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_100 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_99;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_101 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_100;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_102 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_101;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_103 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_102;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_104 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_103;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_105 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_104;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_106 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_105;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_107 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_106;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_108 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_107;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_109 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_108;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_110 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_109;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_111 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_110;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_112 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_111;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_113 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_112;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_114 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_113;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_115 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_114;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_116 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_115;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_117 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_116;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_118 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_117;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_119 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_118;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_120 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_119;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_121 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_120;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_122 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_121;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_123 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_122;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_124 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_123;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_125 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_124;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_126 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_125;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_127 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_126;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_128 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_127;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_129 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_128;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_130 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_129;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_131 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_130;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_132 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_131;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_133 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_132;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_134 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_133;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_135 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_134;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_136 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_135;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_137 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_136;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_138 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_137;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_139 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_138;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_140 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_139;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_141 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_140;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_142 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_141;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_143 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_142;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_144 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_143;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_145 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_144;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_146 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_145;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_147 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_146;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_148 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_147;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_149 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_148;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_150 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_149;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_151 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_150;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_152 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_151;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_153 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_152;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_154 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_153;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_155 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_154;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_156 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_155;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_157 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_156;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_158 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_157;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_159 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_158;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_160 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_159;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_161 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_160;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_162 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_161;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_163 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_162;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_164 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_163;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_165 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_164;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_166 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_165;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_167 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_166;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_168 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_167;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_169 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_168;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_170 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_169;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_171 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_170;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_172 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_171;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_173 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_172;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_174 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_173;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_175 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_174;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_176 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_175;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_177 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_176;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_178 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_177;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_179 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_178;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_180 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_179;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_181 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57_stage_180;
      dark_dark_weights_update_0_read_read_8_stage_14 <= dark_dark_weights_update_0_read_read_8;
      dark_dark_weights_update_0_read_read_8_stage_15 <= dark_dark_weights_update_0_read_read_8_stage_14;
      dark_dark_weights_update_0_read_read_8_stage_16 <= dark_dark_weights_update_0_read_read_8_stage_15;
      dark_dark_weights_update_0_read_read_8_stage_17 <= dark_dark_weights_update_0_read_read_8_stage_16;
      dark_dark_weights_update_0_read_read_8_stage_18 <= dark_dark_weights_update_0_read_read_8_stage_17;
      dark_dark_weights_update_0_read_read_8_stage_19 <= dark_dark_weights_update_0_read_read_8_stage_18;
      dark_dark_weights_update_0_read_read_8_stage_20 <= dark_dark_weights_update_0_read_read_8_stage_19;
      dark_dark_weights_update_0_read_read_8_stage_21 <= dark_dark_weights_update_0_read_read_8_stage_20;
      dark_dark_weights_update_0_read_read_8_stage_22 <= dark_dark_weights_update_0_read_read_8_stage_21;
      dark_dark_weights_update_0_read_read_8_stage_23 <= dark_dark_weights_update_0_read_read_8_stage_22;
      dark_dark_weights_update_0_read_read_8_stage_24 <= dark_dark_weights_update_0_read_read_8_stage_23;
      dark_dark_weights_update_0_read_read_8_stage_25 <= dark_dark_weights_update_0_read_read_8_stage_24;
      dark_dark_weights_update_0_read_read_8_stage_26 <= dark_dark_weights_update_0_read_read_8_stage_25;
      dark_dark_weights_update_0_read_read_8_stage_27 <= dark_dark_weights_update_0_read_read_8_stage_26;
      dark_dark_weights_update_0_read_read_8_stage_28 <= dark_dark_weights_update_0_read_read_8_stage_27;
      dark_dark_weights_update_0_read_read_8_stage_29 <= dark_dark_weights_update_0_read_read_8_stage_28;
      dark_dark_weights_update_0_read_read_8_stage_30 <= dark_dark_weights_update_0_read_read_8_stage_29;
      dark_dark_weights_update_0_read_read_8_stage_31 <= dark_dark_weights_update_0_read_read_8_stage_30;
      dark_dark_weights_update_0_read_read_8_stage_32 <= dark_dark_weights_update_0_read_read_8_stage_31;
      dark_dark_weights_update_0_read_read_8_stage_33 <= dark_dark_weights_update_0_read_read_8_stage_32;
      dark_dark_weights_update_0_read_read_8_stage_34 <= dark_dark_weights_update_0_read_read_8_stage_33;
      dark_dark_weights_update_0_read_read_8_stage_35 <= dark_dark_weights_update_0_read_read_8_stage_34;
      dark_dark_weights_update_0_read_read_8_stage_36 <= dark_dark_weights_update_0_read_read_8_stage_35;
      dark_dark_weights_update_0_read_read_8_stage_37 <= dark_dark_weights_update_0_read_read_8_stage_36;
      dark_dark_weights_update_0_read_read_8_stage_38 <= dark_dark_weights_update_0_read_read_8_stage_37;
      dark_dark_weights_update_0_read_read_8_stage_39 <= dark_dark_weights_update_0_read_read_8_stage_38;
      dark_dark_weights_update_0_read_read_8_stage_40 <= dark_dark_weights_update_0_read_read_8_stage_39;
      dark_dark_weights_update_0_read_read_8_stage_41 <= dark_dark_weights_update_0_read_read_8_stage_40;
      dark_dark_weights_update_0_read_read_8_stage_42 <= dark_dark_weights_update_0_read_read_8_stage_41;
      dark_dark_weights_update_0_read_read_8_stage_43 <= dark_dark_weights_update_0_read_read_8_stage_42;
      dark_dark_weights_update_0_read_read_8_stage_44 <= dark_dark_weights_update_0_read_read_8_stage_43;
      dark_dark_weights_update_0_read_read_8_stage_45 <= dark_dark_weights_update_0_read_read_8_stage_44;
      dark_dark_weights_update_0_read_read_8_stage_46 <= dark_dark_weights_update_0_read_read_8_stage_45;
      dark_dark_weights_update_0_read_read_8_stage_47 <= dark_dark_weights_update_0_read_read_8_stage_46;
      dark_dark_weights_update_0_read_read_8_stage_48 <= dark_dark_weights_update_0_read_read_8_stage_47;
      dark_dark_weights_update_0_read_read_8_stage_49 <= dark_dark_weights_update_0_read_read_8_stage_48;
      dark_dark_weights_update_0_read_read_8_stage_50 <= dark_dark_weights_update_0_read_read_8_stage_49;
      dark_dark_weights_update_0_read_read_8_stage_51 <= dark_dark_weights_update_0_read_read_8_stage_50;
      dark_dark_weights_update_0_read_read_8_stage_52 <= dark_dark_weights_update_0_read_read_8_stage_51;
      dark_dark_weights_update_0_read_read_8_stage_53 <= dark_dark_weights_update_0_read_read_8_stage_52;
      dark_dark_weights_update_0_read_read_8_stage_54 <= dark_dark_weights_update_0_read_read_8_stage_53;
      dark_dark_weights_update_0_read_read_8_stage_55 <= dark_dark_weights_update_0_read_read_8_stage_54;
      dark_dark_weights_update_0_read_read_8_stage_56 <= dark_dark_weights_update_0_read_read_8_stage_55;
      dark_dark_weights_update_0_read_read_8_stage_57 <= dark_dark_weights_update_0_read_read_8_stage_56;
      dark_dark_weights_update_0_read_read_8_stage_58 <= dark_dark_weights_update_0_read_read_8_stage_57;
      dark_dark_weights_update_0_read_read_8_stage_59 <= dark_dark_weights_update_0_read_read_8_stage_58;
      dark_dark_weights_update_0_read_read_8_stage_60 <= dark_dark_weights_update_0_read_read_8_stage_59;
      dark_dark_weights_update_0_read_read_8_stage_61 <= dark_dark_weights_update_0_read_read_8_stage_60;
      dark_dark_weights_update_0_read_read_8_stage_62 <= dark_dark_weights_update_0_read_read_8_stage_61;
      dark_dark_weights_update_0_read_read_8_stage_63 <= dark_dark_weights_update_0_read_read_8_stage_62;
      dark_dark_weights_update_0_read_read_8_stage_64 <= dark_dark_weights_update_0_read_read_8_stage_63;
      dark_dark_weights_update_0_read_read_8_stage_65 <= dark_dark_weights_update_0_read_read_8_stage_64;
      dark_dark_weights_update_0_read_read_8_stage_66 <= dark_dark_weights_update_0_read_read_8_stage_65;
      dark_dark_weights_update_0_read_read_8_stage_67 <= dark_dark_weights_update_0_read_read_8_stage_66;
      dark_dark_weights_update_0_read_read_8_stage_68 <= dark_dark_weights_update_0_read_read_8_stage_67;
      dark_dark_weights_update_0_read_read_8_stage_69 <= dark_dark_weights_update_0_read_read_8_stage_68;
      dark_dark_weights_update_0_read_read_8_stage_70 <= dark_dark_weights_update_0_read_read_8_stage_69;
      dark_dark_weights_update_0_read_read_8_stage_71 <= dark_dark_weights_update_0_read_read_8_stage_70;
      dark_dark_weights_update_0_read_read_8_stage_72 <= dark_dark_weights_update_0_read_read_8_stage_71;
      dark_dark_weights_update_0_read_read_8_stage_73 <= dark_dark_weights_update_0_read_read_8_stage_72;
      dark_dark_weights_update_0_read_read_8_stage_74 <= dark_dark_weights_update_0_read_read_8_stage_73;
      dark_dark_weights_update_0_read_read_8_stage_75 <= dark_dark_weights_update_0_read_read_8_stage_74;
      dark_dark_weights_update_0_read_read_8_stage_76 <= dark_dark_weights_update_0_read_read_8_stage_75;
      dark_dark_weights_update_0_read_read_8_stage_77 <= dark_dark_weights_update_0_read_read_8_stage_76;
      dark_dark_weights_update_0_read_read_8_stage_78 <= dark_dark_weights_update_0_read_read_8_stage_77;
      dark_dark_weights_update_0_read_read_8_stage_79 <= dark_dark_weights_update_0_read_read_8_stage_78;
      dark_dark_weights_update_0_read_read_8_stage_80 <= dark_dark_weights_update_0_read_read_8_stage_79;
      dark_dark_weights_update_0_read_read_8_stage_81 <= dark_dark_weights_update_0_read_read_8_stage_80;
      dark_dark_weights_update_0_read_read_8_stage_82 <= dark_dark_weights_update_0_read_read_8_stage_81;
      dark_dark_weights_update_0_read_read_8_stage_83 <= dark_dark_weights_update_0_read_read_8_stage_82;
      dark_dark_weights_update_0_read_read_8_stage_84 <= dark_dark_weights_update_0_read_read_8_stage_83;
      dark_dark_weights_update_0_read_read_8_stage_85 <= dark_dark_weights_update_0_read_read_8_stage_84;
      dark_dark_weights_update_0_read_read_8_stage_86 <= dark_dark_weights_update_0_read_read_8_stage_85;
      dark_dark_weights_update_0_read_read_8_stage_87 <= dark_dark_weights_update_0_read_read_8_stage_86;
      dark_dark_weights_update_0_read_read_8_stage_88 <= dark_dark_weights_update_0_read_read_8_stage_87;
      dark_dark_weights_update_0_read_read_8_stage_89 <= dark_dark_weights_update_0_read_read_8_stage_88;
      dark_dark_weights_update_0_read_read_8_stage_90 <= dark_dark_weights_update_0_read_read_8_stage_89;
      dark_dark_weights_update_0_read_read_8_stage_91 <= dark_dark_weights_update_0_read_read_8_stage_90;
      dark_dark_weights_update_0_read_read_8_stage_92 <= dark_dark_weights_update_0_read_read_8_stage_91;
      dark_dark_weights_update_0_read_read_8_stage_93 <= dark_dark_weights_update_0_read_read_8_stage_92;
      dark_dark_weights_update_0_read_read_8_stage_94 <= dark_dark_weights_update_0_read_read_8_stage_93;
      dark_dark_weights_update_0_read_read_8_stage_95 <= dark_dark_weights_update_0_read_read_8_stage_94;
      dark_dark_weights_update_0_read_read_8_stage_96 <= dark_dark_weights_update_0_read_read_8_stage_95;
      dark_dark_weights_update_0_read_read_8_stage_97 <= dark_dark_weights_update_0_read_read_8_stage_96;
      dark_dark_weights_update_0_read_read_8_stage_98 <= dark_dark_weights_update_0_read_read_8_stage_97;
      dark_dark_weights_update_0_read_read_8_stage_99 <= dark_dark_weights_update_0_read_read_8_stage_98;
      dark_dark_weights_update_0_read_read_8_stage_100 <= dark_dark_weights_update_0_read_read_8_stage_99;
      dark_dark_weights_update_0_read_read_8_stage_101 <= dark_dark_weights_update_0_read_read_8_stage_100;
      dark_dark_weights_update_0_read_read_8_stage_102 <= dark_dark_weights_update_0_read_read_8_stage_101;
      dark_dark_weights_update_0_read_read_8_stage_103 <= dark_dark_weights_update_0_read_read_8_stage_102;
      dark_dark_weights_update_0_read_read_8_stage_104 <= dark_dark_weights_update_0_read_read_8_stage_103;
      dark_dark_weights_update_0_read_read_8_stage_105 <= dark_dark_weights_update_0_read_read_8_stage_104;
      dark_dark_weights_update_0_read_read_8_stage_106 <= dark_dark_weights_update_0_read_read_8_stage_105;
      dark_dark_weights_update_0_read_read_8_stage_107 <= dark_dark_weights_update_0_read_read_8_stage_106;
      dark_dark_weights_update_0_read_read_8_stage_108 <= dark_dark_weights_update_0_read_read_8_stage_107;
      dark_dark_weights_update_0_read_read_8_stage_109 <= dark_dark_weights_update_0_read_read_8_stage_108;
      dark_dark_weights_update_0_read_read_8_stage_110 <= dark_dark_weights_update_0_read_read_8_stage_109;
      dark_dark_weights_update_0_read_read_8_stage_111 <= dark_dark_weights_update_0_read_read_8_stage_110;
      dark_dark_weights_update_0_read_read_8_stage_112 <= dark_dark_weights_update_0_read_read_8_stage_111;
      dark_dark_weights_update_0_read_read_8_stage_113 <= dark_dark_weights_update_0_read_read_8_stage_112;
      dark_dark_weights_update_0_read_read_8_stage_114 <= dark_dark_weights_update_0_read_read_8_stage_113;
      dark_dark_weights_update_0_read_read_8_stage_115 <= dark_dark_weights_update_0_read_read_8_stage_114;
      dark_dark_weights_update_0_read_read_8_stage_116 <= dark_dark_weights_update_0_read_read_8_stage_115;
      dark_dark_weights_update_0_read_read_8_stage_117 <= dark_dark_weights_update_0_read_read_8_stage_116;
      dark_dark_weights_update_0_read_read_8_stage_118 <= dark_dark_weights_update_0_read_read_8_stage_117;
      dark_dark_weights_update_0_read_read_8_stage_119 <= dark_dark_weights_update_0_read_read_8_stage_118;
      dark_dark_weights_update_0_read_read_8_stage_120 <= dark_dark_weights_update_0_read_read_8_stage_119;
      dark_dark_weights_update_0_read_read_8_stage_121 <= dark_dark_weights_update_0_read_read_8_stage_120;
      dark_dark_weights_update_0_read_read_8_stage_122 <= dark_dark_weights_update_0_read_read_8_stage_121;
      dark_dark_weights_update_0_read_read_8_stage_123 <= dark_dark_weights_update_0_read_read_8_stage_122;
      dark_dark_weights_update_0_read_read_8_stage_124 <= dark_dark_weights_update_0_read_read_8_stage_123;
      dark_dark_weights_update_0_read_read_8_stage_125 <= dark_dark_weights_update_0_read_read_8_stage_124;
      dark_dark_weights_update_0_read_read_8_stage_126 <= dark_dark_weights_update_0_read_read_8_stage_125;
      dark_dark_weights_update_0_read_read_8_stage_127 <= dark_dark_weights_update_0_read_read_8_stage_126;
      dark_dark_weights_update_0_read_read_8_stage_128 <= dark_dark_weights_update_0_read_read_8_stage_127;
      dark_dark_weights_update_0_read_read_8_stage_129 <= dark_dark_weights_update_0_read_read_8_stage_128;
      dark_dark_weights_update_0_read_read_8_stage_130 <= dark_dark_weights_update_0_read_read_8_stage_129;
      dark_dark_weights_update_0_read_read_8_stage_131 <= dark_dark_weights_update_0_read_read_8_stage_130;
      dark_dark_weights_update_0_read_read_8_stage_132 <= dark_dark_weights_update_0_read_read_8_stage_131;
      dark_dark_weights_update_0_read_read_8_stage_133 <= dark_dark_weights_update_0_read_read_8_stage_132;
      dark_dark_weights_update_0_read_read_8_stage_134 <= dark_dark_weights_update_0_read_read_8_stage_133;
      dark_dark_weights_update_0_read_read_8_stage_135 <= dark_dark_weights_update_0_read_read_8_stage_134;
      dark_dark_weights_update_0_read_read_8_stage_136 <= dark_dark_weights_update_0_read_read_8_stage_135;
      dark_dark_weights_update_0_read_read_8_stage_137 <= dark_dark_weights_update_0_read_read_8_stage_136;
      dark_dark_weights_update_0_read_read_8_stage_138 <= dark_dark_weights_update_0_read_read_8_stage_137;
      dark_dark_weights_update_0_read_read_8_stage_139 <= dark_dark_weights_update_0_read_read_8_stage_138;
      dark_dark_weights_update_0_read_read_8_stage_140 <= dark_dark_weights_update_0_read_read_8_stage_139;
      dark_dark_weights_update_0_read_read_8_stage_141 <= dark_dark_weights_update_0_read_read_8_stage_140;
      dark_dark_weights_update_0_read_read_8_stage_142 <= dark_dark_weights_update_0_read_read_8_stage_141;
      dark_dark_weights_update_0_read_read_8_stage_143 <= dark_dark_weights_update_0_read_read_8_stage_142;
      dark_dark_weights_update_0_read_read_8_stage_144 <= dark_dark_weights_update_0_read_read_8_stage_143;
      dark_dark_weights_update_0_read_read_8_stage_145 <= dark_dark_weights_update_0_read_read_8_stage_144;
      dark_dark_weights_update_0_read_read_8_stage_146 <= dark_dark_weights_update_0_read_read_8_stage_145;
      dark_dark_weights_update_0_read_read_8_stage_147 <= dark_dark_weights_update_0_read_read_8_stage_146;
      dark_dark_weights_update_0_read_read_8_stage_148 <= dark_dark_weights_update_0_read_read_8_stage_147;
      dark_dark_weights_update_0_read_read_8_stage_149 <= dark_dark_weights_update_0_read_read_8_stage_148;
      dark_dark_weights_update_0_read_read_8_stage_150 <= dark_dark_weights_update_0_read_read_8_stage_149;
      dark_dark_weights_update_0_read_read_8_stage_151 <= dark_dark_weights_update_0_read_read_8_stage_150;
      dark_dark_weights_update_0_read_read_8_stage_152 <= dark_dark_weights_update_0_read_read_8_stage_151;
      dark_dark_weights_update_0_read_read_8_stage_153 <= dark_dark_weights_update_0_read_read_8_stage_152;
      dark_dark_weights_update_0_read_read_8_stage_154 <= dark_dark_weights_update_0_read_read_8_stage_153;
      dark_dark_weights_update_0_read_read_8_stage_155 <= dark_dark_weights_update_0_read_read_8_stage_154;
      dark_dark_weights_update_0_read_read_8_stage_156 <= dark_dark_weights_update_0_read_read_8_stage_155;
      dark_dark_weights_update_0_read_read_8_stage_157 <= dark_dark_weights_update_0_read_read_8_stage_156;
      dark_dark_weights_update_0_read_read_8_stage_158 <= dark_dark_weights_update_0_read_read_8_stage_157;
      dark_dark_weights_update_0_read_read_8_stage_159 <= dark_dark_weights_update_0_read_read_8_stage_158;
      dark_dark_weights_update_0_read_read_8_stage_160 <= dark_dark_weights_update_0_read_read_8_stage_159;
      dark_dark_weights_update_0_read_read_8_stage_161 <= dark_dark_weights_update_0_read_read_8_stage_160;
      dark_dark_weights_update_0_read_read_8_stage_162 <= dark_dark_weights_update_0_read_read_8_stage_161;
      dark_dark_weights_update_0_read_read_8_stage_163 <= dark_dark_weights_update_0_read_read_8_stage_162;
      dark_dark_weights_update_0_read_read_8_stage_164 <= dark_dark_weights_update_0_read_read_8_stage_163;
      dark_dark_weights_update_0_read_read_8_stage_165 <= dark_dark_weights_update_0_read_read_8_stage_164;
      dark_dark_weights_update_0_read_read_8_stage_166 <= dark_dark_weights_update_0_read_read_8_stage_165;
      dark_dark_weights_update_0_read_read_8_stage_167 <= dark_dark_weights_update_0_read_read_8_stage_166;
      dark_dark_weights_update_0_read_read_8_stage_168 <= dark_dark_weights_update_0_read_read_8_stage_167;
      dark_dark_weights_update_0_read_read_8_stage_169 <= dark_dark_weights_update_0_read_read_8_stage_168;
      dark_dark_weights_update_0_read_read_8_stage_170 <= dark_dark_weights_update_0_read_read_8_stage_169;
      dark_dark_weights_update_0_read_read_8_stage_171 <= dark_dark_weights_update_0_read_read_8_stage_170;
      dark_dark_weights_update_0_read_read_8_stage_172 <= dark_dark_weights_update_0_read_read_8_stage_171;
      dark_dark_weights_update_0_read_read_8_stage_173 <= dark_dark_weights_update_0_read_read_8_stage_172;
      dark_dark_weights_update_0_read_read_8_stage_174 <= dark_dark_weights_update_0_read_read_8_stage_173;
      dark_dark_weights_update_0_read_read_8_stage_175 <= dark_dark_weights_update_0_read_read_8_stage_174;
      dark_dark_weights_update_0_read_read_8_stage_176 <= dark_dark_weights_update_0_read_read_8_stage_175;
      dark_dark_weights_update_0_read_read_8_stage_177 <= dark_dark_weights_update_0_read_read_8_stage_176;
      dark_dark_weights_update_0_read_read_8_stage_178 <= dark_dark_weights_update_0_read_read_8_stage_177;
      dark_dark_weights_update_0_read_read_8_stage_179 <= dark_dark_weights_update_0_read_read_8_stage_178;
      dark_dark_weights_update_0_read_read_8_stage_180 <= dark_dark_weights_update_0_read_read_8_stage_179;
      dark_dark_weights_update_0_read_read_8_stage_181 <= dark_dark_weights_update_0_read_read_8_stage_180;
      dark_weights_update_0_stage_15 <= dark_weights_update_0;
      dark_weights_update_0_stage_16 <= dark_weights_update_0_stage_15;
      dark_weights_update_0_stage_17 <= dark_weights_update_0_stage_16;
      dark_weights_update_0_stage_18 <= dark_weights_update_0_stage_17;
      dark_weights_update_0_stage_19 <= dark_weights_update_0_stage_18;
      dark_weights_update_0_stage_20 <= dark_weights_update_0_stage_19;
      dark_weights_update_0_stage_21 <= dark_weights_update_0_stage_20;
      dark_weights_update_0_stage_22 <= dark_weights_update_0_stage_21;
      dark_weights_update_0_stage_23 <= dark_weights_update_0_stage_22;
      dark_weights_update_0_stage_24 <= dark_weights_update_0_stage_23;
      dark_weights_update_0_stage_25 <= dark_weights_update_0_stage_24;
      dark_weights_update_0_stage_26 <= dark_weights_update_0_stage_25;
      dark_weights_update_0_stage_27 <= dark_weights_update_0_stage_26;
      dark_weights_update_0_stage_28 <= dark_weights_update_0_stage_27;
      dark_weights_update_0_stage_29 <= dark_weights_update_0_stage_28;
      dark_weights_update_0_stage_30 <= dark_weights_update_0_stage_29;
      dark_weights_update_0_stage_31 <= dark_weights_update_0_stage_30;
      dark_weights_update_0_stage_32 <= dark_weights_update_0_stage_31;
      dark_weights_update_0_stage_33 <= dark_weights_update_0_stage_32;
      dark_weights_update_0_stage_34 <= dark_weights_update_0_stage_33;
      dark_weights_update_0_stage_35 <= dark_weights_update_0_stage_34;
      dark_weights_update_0_stage_36 <= dark_weights_update_0_stage_35;
      dark_weights_update_0_stage_37 <= dark_weights_update_0_stage_36;
      dark_weights_update_0_stage_38 <= dark_weights_update_0_stage_37;
      dark_weights_update_0_stage_39 <= dark_weights_update_0_stage_38;
      dark_weights_update_0_stage_40 <= dark_weights_update_0_stage_39;
      dark_weights_update_0_stage_41 <= dark_weights_update_0_stage_40;
      dark_weights_update_0_stage_42 <= dark_weights_update_0_stage_41;
      dark_weights_update_0_stage_43 <= dark_weights_update_0_stage_42;
      dark_weights_update_0_stage_44 <= dark_weights_update_0_stage_43;
      dark_weights_update_0_stage_45 <= dark_weights_update_0_stage_44;
      dark_weights_update_0_stage_46 <= dark_weights_update_0_stage_45;
      dark_weights_update_0_stage_47 <= dark_weights_update_0_stage_46;
      dark_weights_update_0_stage_48 <= dark_weights_update_0_stage_47;
      dark_weights_update_0_stage_49 <= dark_weights_update_0_stage_48;
      dark_weights_update_0_stage_50 <= dark_weights_update_0_stage_49;
      dark_weights_update_0_stage_51 <= dark_weights_update_0_stage_50;
      dark_weights_update_0_stage_52 <= dark_weights_update_0_stage_51;
      dark_weights_update_0_stage_53 <= dark_weights_update_0_stage_52;
      dark_weights_update_0_stage_54 <= dark_weights_update_0_stage_53;
      dark_weights_update_0_stage_55 <= dark_weights_update_0_stage_54;
      dark_weights_update_0_stage_56 <= dark_weights_update_0_stage_55;
      dark_weights_update_0_stage_57 <= dark_weights_update_0_stage_56;
      dark_weights_update_0_stage_58 <= dark_weights_update_0_stage_57;
      dark_weights_update_0_stage_59 <= dark_weights_update_0_stage_58;
      dark_weights_update_0_stage_60 <= dark_weights_update_0_stage_59;
      dark_weights_update_0_stage_61 <= dark_weights_update_0_stage_60;
      dark_weights_update_0_stage_62 <= dark_weights_update_0_stage_61;
      dark_weights_update_0_stage_63 <= dark_weights_update_0_stage_62;
      dark_weights_update_0_stage_64 <= dark_weights_update_0_stage_63;
      dark_weights_update_0_stage_65 <= dark_weights_update_0_stage_64;
      dark_weights_update_0_stage_66 <= dark_weights_update_0_stage_65;
      dark_weights_update_0_stage_67 <= dark_weights_update_0_stage_66;
      dark_weights_update_0_stage_68 <= dark_weights_update_0_stage_67;
      dark_weights_update_0_stage_69 <= dark_weights_update_0_stage_68;
      dark_weights_update_0_stage_70 <= dark_weights_update_0_stage_69;
      dark_weights_update_0_stage_71 <= dark_weights_update_0_stage_70;
      dark_weights_update_0_stage_72 <= dark_weights_update_0_stage_71;
      dark_weights_update_0_stage_73 <= dark_weights_update_0_stage_72;
      dark_weights_update_0_stage_74 <= dark_weights_update_0_stage_73;
      dark_weights_update_0_stage_75 <= dark_weights_update_0_stage_74;
      dark_weights_update_0_stage_76 <= dark_weights_update_0_stage_75;
      dark_weights_update_0_stage_77 <= dark_weights_update_0_stage_76;
      dark_weights_update_0_stage_78 <= dark_weights_update_0_stage_77;
      dark_weights_update_0_stage_79 <= dark_weights_update_0_stage_78;
      dark_weights_update_0_stage_80 <= dark_weights_update_0_stage_79;
      dark_weights_update_0_stage_81 <= dark_weights_update_0_stage_80;
      dark_weights_update_0_stage_82 <= dark_weights_update_0_stage_81;
      dark_weights_update_0_stage_83 <= dark_weights_update_0_stage_82;
      dark_weights_update_0_stage_84 <= dark_weights_update_0_stage_83;
      dark_weights_update_0_stage_85 <= dark_weights_update_0_stage_84;
      dark_weights_update_0_stage_86 <= dark_weights_update_0_stage_85;
      dark_weights_update_0_stage_87 <= dark_weights_update_0_stage_86;
      dark_weights_update_0_stage_88 <= dark_weights_update_0_stage_87;
      dark_weights_update_0_stage_89 <= dark_weights_update_0_stage_88;
      dark_weights_update_0_stage_90 <= dark_weights_update_0_stage_89;
      dark_weights_update_0_stage_91 <= dark_weights_update_0_stage_90;
      dark_weights_update_0_stage_92 <= dark_weights_update_0_stage_91;
      dark_weights_update_0_stage_93 <= dark_weights_update_0_stage_92;
      dark_weights_update_0_stage_94 <= dark_weights_update_0_stage_93;
      dark_weights_update_0_stage_95 <= dark_weights_update_0_stage_94;
      dark_weights_update_0_stage_96 <= dark_weights_update_0_stage_95;
      dark_weights_update_0_stage_97 <= dark_weights_update_0_stage_96;
      dark_weights_update_0_stage_98 <= dark_weights_update_0_stage_97;
      dark_weights_update_0_stage_99 <= dark_weights_update_0_stage_98;
      dark_weights_update_0_stage_100 <= dark_weights_update_0_stage_99;
      dark_weights_update_0_stage_101 <= dark_weights_update_0_stage_100;
      dark_weights_update_0_stage_102 <= dark_weights_update_0_stage_101;
      dark_weights_update_0_stage_103 <= dark_weights_update_0_stage_102;
      dark_weights_update_0_stage_104 <= dark_weights_update_0_stage_103;
      dark_weights_update_0_stage_105 <= dark_weights_update_0_stage_104;
      dark_weights_update_0_stage_106 <= dark_weights_update_0_stage_105;
      dark_weights_update_0_stage_107 <= dark_weights_update_0_stage_106;
      dark_weights_update_0_stage_108 <= dark_weights_update_0_stage_107;
      dark_weights_update_0_stage_109 <= dark_weights_update_0_stage_108;
      dark_weights_update_0_stage_110 <= dark_weights_update_0_stage_109;
      dark_weights_update_0_stage_111 <= dark_weights_update_0_stage_110;
      dark_weights_update_0_stage_112 <= dark_weights_update_0_stage_111;
      dark_weights_update_0_stage_113 <= dark_weights_update_0_stage_112;
      dark_weights_update_0_stage_114 <= dark_weights_update_0_stage_113;
      dark_weights_update_0_stage_115 <= dark_weights_update_0_stage_114;
      dark_weights_update_0_stage_116 <= dark_weights_update_0_stage_115;
      dark_weights_update_0_stage_117 <= dark_weights_update_0_stage_116;
      dark_weights_update_0_stage_118 <= dark_weights_update_0_stage_117;
      dark_weights_update_0_stage_119 <= dark_weights_update_0_stage_118;
      dark_weights_update_0_stage_120 <= dark_weights_update_0_stage_119;
      dark_weights_update_0_stage_121 <= dark_weights_update_0_stage_120;
      dark_weights_update_0_stage_122 <= dark_weights_update_0_stage_121;
      dark_weights_update_0_stage_123 <= dark_weights_update_0_stage_122;
      dark_weights_update_0_stage_124 <= dark_weights_update_0_stage_123;
      dark_weights_update_0_stage_125 <= dark_weights_update_0_stage_124;
      dark_weights_update_0_stage_126 <= dark_weights_update_0_stage_125;
      dark_weights_update_0_stage_127 <= dark_weights_update_0_stage_126;
      dark_weights_update_0_stage_128 <= dark_weights_update_0_stage_127;
      dark_weights_update_0_stage_129 <= dark_weights_update_0_stage_128;
      dark_weights_update_0_stage_130 <= dark_weights_update_0_stage_129;
      dark_weights_update_0_stage_131 <= dark_weights_update_0_stage_130;
      dark_weights_update_0_stage_132 <= dark_weights_update_0_stage_131;
      dark_weights_update_0_stage_133 <= dark_weights_update_0_stage_132;
      dark_weights_update_0_stage_134 <= dark_weights_update_0_stage_133;
      dark_weights_update_0_stage_135 <= dark_weights_update_0_stage_134;
      dark_weights_update_0_stage_136 <= dark_weights_update_0_stage_135;
      dark_weights_update_0_stage_137 <= dark_weights_update_0_stage_136;
      dark_weights_update_0_stage_138 <= dark_weights_update_0_stage_137;
      dark_weights_update_0_stage_139 <= dark_weights_update_0_stage_138;
      dark_weights_update_0_stage_140 <= dark_weights_update_0_stage_139;
      dark_weights_update_0_stage_141 <= dark_weights_update_0_stage_140;
      dark_weights_update_0_stage_142 <= dark_weights_update_0_stage_141;
      dark_weights_update_0_stage_143 <= dark_weights_update_0_stage_142;
      dark_weights_update_0_stage_144 <= dark_weights_update_0_stage_143;
      dark_weights_update_0_stage_145 <= dark_weights_update_0_stage_144;
      dark_weights_update_0_stage_146 <= dark_weights_update_0_stage_145;
      dark_weights_update_0_stage_147 <= dark_weights_update_0_stage_146;
      dark_weights_update_0_stage_148 <= dark_weights_update_0_stage_147;
      dark_weights_update_0_stage_149 <= dark_weights_update_0_stage_148;
      dark_weights_update_0_stage_150 <= dark_weights_update_0_stage_149;
      dark_weights_update_0_stage_151 <= dark_weights_update_0_stage_150;
      dark_weights_update_0_stage_152 <= dark_weights_update_0_stage_151;
      dark_weights_update_0_stage_153 <= dark_weights_update_0_stage_152;
      dark_weights_update_0_stage_154 <= dark_weights_update_0_stage_153;
      dark_weights_update_0_stage_155 <= dark_weights_update_0_stage_154;
      dark_weights_update_0_stage_156 <= dark_weights_update_0_stage_155;
      dark_weights_update_0_stage_157 <= dark_weights_update_0_stage_156;
      dark_weights_update_0_stage_158 <= dark_weights_update_0_stage_157;
      dark_weights_update_0_stage_159 <= dark_weights_update_0_stage_158;
      dark_weights_update_0_stage_160 <= dark_weights_update_0_stage_159;
      dark_weights_update_0_stage_161 <= dark_weights_update_0_stage_160;
      dark_weights_update_0_stage_162 <= dark_weights_update_0_stage_161;
      dark_weights_update_0_stage_163 <= dark_weights_update_0_stage_162;
      dark_weights_update_0_stage_164 <= dark_weights_update_0_stage_163;
      dark_weights_update_0_stage_165 <= dark_weights_update_0_stage_164;
      dark_weights_update_0_stage_166 <= dark_weights_update_0_stage_165;
      dark_weights_update_0_stage_167 <= dark_weights_update_0_stage_166;
      dark_weights_update_0_stage_168 <= dark_weights_update_0_stage_167;
      dark_weights_update_0_stage_169 <= dark_weights_update_0_stage_168;
      dark_weights_update_0_stage_170 <= dark_weights_update_0_stage_169;
      dark_weights_update_0_stage_171 <= dark_weights_update_0_stage_170;
      dark_weights_update_0_stage_172 <= dark_weights_update_0_stage_171;
      dark_weights_update_0_stage_173 <= dark_weights_update_0_stage_172;
      dark_weights_update_0_stage_174 <= dark_weights_update_0_stage_173;
      dark_weights_update_0_stage_175 <= dark_weights_update_0_stage_174;
      dark_weights_update_0_stage_176 <= dark_weights_update_0_stage_175;
      dark_weights_update_0_stage_177 <= dark_weights_update_0_stage_176;
      dark_weights_update_0_stage_178 <= dark_weights_update_0_stage_177;
      dark_weights_update_0_stage_179 <= dark_weights_update_0_stage_178;
      dark_weights_update_0_stage_180 <= dark_weights_update_0_stage_179;
      dark_weights_update_0_stage_181 <= dark_weights_update_0_stage_180;
      dark_weights_dark_weights_update_0_write_write_9_stage_16 <= dark_weights_dark_weights_update_0_write_write_9;
      dark_weights_dark_weights_update_0_write_write_9_stage_17 <= dark_weights_dark_weights_update_0_write_write_9_stage_16;
      dark_weights_dark_weights_update_0_write_write_9_stage_18 <= dark_weights_dark_weights_update_0_write_write_9_stage_17;
      dark_weights_dark_weights_update_0_write_write_9_stage_19 <= dark_weights_dark_weights_update_0_write_write_9_stage_18;
      dark_weights_dark_weights_update_0_write_write_9_stage_20 <= dark_weights_dark_weights_update_0_write_write_9_stage_19;
      dark_weights_dark_weights_update_0_write_write_9_stage_21 <= dark_weights_dark_weights_update_0_write_write_9_stage_20;
      dark_weights_dark_weights_update_0_write_write_9_stage_22 <= dark_weights_dark_weights_update_0_write_write_9_stage_21;
      dark_weights_dark_weights_update_0_write_write_9_stage_23 <= dark_weights_dark_weights_update_0_write_write_9_stage_22;
      dark_weights_dark_weights_update_0_write_write_9_stage_24 <= dark_weights_dark_weights_update_0_write_write_9_stage_23;
      dark_weights_dark_weights_update_0_write_write_9_stage_25 <= dark_weights_dark_weights_update_0_write_write_9_stage_24;
      dark_weights_dark_weights_update_0_write_write_9_stage_26 <= dark_weights_dark_weights_update_0_write_write_9_stage_25;
      dark_weights_dark_weights_update_0_write_write_9_stage_27 <= dark_weights_dark_weights_update_0_write_write_9_stage_26;
      dark_weights_dark_weights_update_0_write_write_9_stage_28 <= dark_weights_dark_weights_update_0_write_write_9_stage_27;
      dark_weights_dark_weights_update_0_write_write_9_stage_29 <= dark_weights_dark_weights_update_0_write_write_9_stage_28;
      dark_weights_dark_weights_update_0_write_write_9_stage_30 <= dark_weights_dark_weights_update_0_write_write_9_stage_29;
      dark_weights_dark_weights_update_0_write_write_9_stage_31 <= dark_weights_dark_weights_update_0_write_write_9_stage_30;
      dark_weights_dark_weights_update_0_write_write_9_stage_32 <= dark_weights_dark_weights_update_0_write_write_9_stage_31;
      dark_weights_dark_weights_update_0_write_write_9_stage_33 <= dark_weights_dark_weights_update_0_write_write_9_stage_32;
      dark_weights_dark_weights_update_0_write_write_9_stage_34 <= dark_weights_dark_weights_update_0_write_write_9_stage_33;
      dark_weights_dark_weights_update_0_write_write_9_stage_35 <= dark_weights_dark_weights_update_0_write_write_9_stage_34;
      dark_weights_dark_weights_update_0_write_write_9_stage_36 <= dark_weights_dark_weights_update_0_write_write_9_stage_35;
      dark_weights_dark_weights_update_0_write_write_9_stage_37 <= dark_weights_dark_weights_update_0_write_write_9_stage_36;
      dark_weights_dark_weights_update_0_write_write_9_stage_38 <= dark_weights_dark_weights_update_0_write_write_9_stage_37;
      dark_weights_dark_weights_update_0_write_write_9_stage_39 <= dark_weights_dark_weights_update_0_write_write_9_stage_38;
      dark_weights_dark_weights_update_0_write_write_9_stage_40 <= dark_weights_dark_weights_update_0_write_write_9_stage_39;
      dark_weights_dark_weights_update_0_write_write_9_stage_41 <= dark_weights_dark_weights_update_0_write_write_9_stage_40;
      dark_weights_dark_weights_update_0_write_write_9_stage_42 <= dark_weights_dark_weights_update_0_write_write_9_stage_41;
      dark_weights_dark_weights_update_0_write_write_9_stage_43 <= dark_weights_dark_weights_update_0_write_write_9_stage_42;
      dark_weights_dark_weights_update_0_write_write_9_stage_44 <= dark_weights_dark_weights_update_0_write_write_9_stage_43;
      dark_weights_dark_weights_update_0_write_write_9_stage_45 <= dark_weights_dark_weights_update_0_write_write_9_stage_44;
      dark_weights_dark_weights_update_0_write_write_9_stage_46 <= dark_weights_dark_weights_update_0_write_write_9_stage_45;
      dark_weights_dark_weights_update_0_write_write_9_stage_47 <= dark_weights_dark_weights_update_0_write_write_9_stage_46;
      dark_weights_dark_weights_update_0_write_write_9_stage_48 <= dark_weights_dark_weights_update_0_write_write_9_stage_47;
      dark_weights_dark_weights_update_0_write_write_9_stage_49 <= dark_weights_dark_weights_update_0_write_write_9_stage_48;
      dark_weights_dark_weights_update_0_write_write_9_stage_50 <= dark_weights_dark_weights_update_0_write_write_9_stage_49;
      dark_weights_dark_weights_update_0_write_write_9_stage_51 <= dark_weights_dark_weights_update_0_write_write_9_stage_50;
      dark_weights_dark_weights_update_0_write_write_9_stage_52 <= dark_weights_dark_weights_update_0_write_write_9_stage_51;
      dark_weights_dark_weights_update_0_write_write_9_stage_53 <= dark_weights_dark_weights_update_0_write_write_9_stage_52;
      dark_weights_dark_weights_update_0_write_write_9_stage_54 <= dark_weights_dark_weights_update_0_write_write_9_stage_53;
      dark_weights_dark_weights_update_0_write_write_9_stage_55 <= dark_weights_dark_weights_update_0_write_write_9_stage_54;
      dark_weights_dark_weights_update_0_write_write_9_stage_56 <= dark_weights_dark_weights_update_0_write_write_9_stage_55;
      dark_weights_dark_weights_update_0_write_write_9_stage_57 <= dark_weights_dark_weights_update_0_write_write_9_stage_56;
      dark_weights_dark_weights_update_0_write_write_9_stage_58 <= dark_weights_dark_weights_update_0_write_write_9_stage_57;
      dark_weights_dark_weights_update_0_write_write_9_stage_59 <= dark_weights_dark_weights_update_0_write_write_9_stage_58;
      dark_weights_dark_weights_update_0_write_write_9_stage_60 <= dark_weights_dark_weights_update_0_write_write_9_stage_59;
      dark_weights_dark_weights_update_0_write_write_9_stage_61 <= dark_weights_dark_weights_update_0_write_write_9_stage_60;
      dark_weights_dark_weights_update_0_write_write_9_stage_62 <= dark_weights_dark_weights_update_0_write_write_9_stage_61;
      dark_weights_dark_weights_update_0_write_write_9_stage_63 <= dark_weights_dark_weights_update_0_write_write_9_stage_62;
      dark_weights_dark_weights_update_0_write_write_9_stage_64 <= dark_weights_dark_weights_update_0_write_write_9_stage_63;
      dark_weights_dark_weights_update_0_write_write_9_stage_65 <= dark_weights_dark_weights_update_0_write_write_9_stage_64;
      dark_weights_dark_weights_update_0_write_write_9_stage_66 <= dark_weights_dark_weights_update_0_write_write_9_stage_65;
      dark_weights_dark_weights_update_0_write_write_9_stage_67 <= dark_weights_dark_weights_update_0_write_write_9_stage_66;
      dark_weights_dark_weights_update_0_write_write_9_stage_68 <= dark_weights_dark_weights_update_0_write_write_9_stage_67;
      dark_weights_dark_weights_update_0_write_write_9_stage_69 <= dark_weights_dark_weights_update_0_write_write_9_stage_68;
      dark_weights_dark_weights_update_0_write_write_9_stage_70 <= dark_weights_dark_weights_update_0_write_write_9_stage_69;
      dark_weights_dark_weights_update_0_write_write_9_stage_71 <= dark_weights_dark_weights_update_0_write_write_9_stage_70;
      dark_weights_dark_weights_update_0_write_write_9_stage_72 <= dark_weights_dark_weights_update_0_write_write_9_stage_71;
      dark_weights_dark_weights_update_0_write_write_9_stage_73 <= dark_weights_dark_weights_update_0_write_write_9_stage_72;
      dark_weights_dark_weights_update_0_write_write_9_stage_74 <= dark_weights_dark_weights_update_0_write_write_9_stage_73;
      dark_weights_dark_weights_update_0_write_write_9_stage_75 <= dark_weights_dark_weights_update_0_write_write_9_stage_74;
      dark_weights_dark_weights_update_0_write_write_9_stage_76 <= dark_weights_dark_weights_update_0_write_write_9_stage_75;
      dark_weights_dark_weights_update_0_write_write_9_stage_77 <= dark_weights_dark_weights_update_0_write_write_9_stage_76;
      dark_weights_dark_weights_update_0_write_write_9_stage_78 <= dark_weights_dark_weights_update_0_write_write_9_stage_77;
      dark_weights_dark_weights_update_0_write_write_9_stage_79 <= dark_weights_dark_weights_update_0_write_write_9_stage_78;
      dark_weights_dark_weights_update_0_write_write_9_stage_80 <= dark_weights_dark_weights_update_0_write_write_9_stage_79;
      dark_weights_dark_weights_update_0_write_write_9_stage_81 <= dark_weights_dark_weights_update_0_write_write_9_stage_80;
      dark_weights_dark_weights_update_0_write_write_9_stage_82 <= dark_weights_dark_weights_update_0_write_write_9_stage_81;
      dark_weights_dark_weights_update_0_write_write_9_stage_83 <= dark_weights_dark_weights_update_0_write_write_9_stage_82;
      dark_weights_dark_weights_update_0_write_write_9_stage_84 <= dark_weights_dark_weights_update_0_write_write_9_stage_83;
      dark_weights_dark_weights_update_0_write_write_9_stage_85 <= dark_weights_dark_weights_update_0_write_write_9_stage_84;
      dark_weights_dark_weights_update_0_write_write_9_stage_86 <= dark_weights_dark_weights_update_0_write_write_9_stage_85;
      dark_weights_dark_weights_update_0_write_write_9_stage_87 <= dark_weights_dark_weights_update_0_write_write_9_stage_86;
      dark_weights_dark_weights_update_0_write_write_9_stage_88 <= dark_weights_dark_weights_update_0_write_write_9_stage_87;
      dark_weights_dark_weights_update_0_write_write_9_stage_89 <= dark_weights_dark_weights_update_0_write_write_9_stage_88;
      dark_weights_dark_weights_update_0_write_write_9_stage_90 <= dark_weights_dark_weights_update_0_write_write_9_stage_89;
      dark_weights_dark_weights_update_0_write_write_9_stage_91 <= dark_weights_dark_weights_update_0_write_write_9_stage_90;
      dark_weights_dark_weights_update_0_write_write_9_stage_92 <= dark_weights_dark_weights_update_0_write_write_9_stage_91;
      dark_weights_dark_weights_update_0_write_write_9_stage_93 <= dark_weights_dark_weights_update_0_write_write_9_stage_92;
      dark_weights_dark_weights_update_0_write_write_9_stage_94 <= dark_weights_dark_weights_update_0_write_write_9_stage_93;
      dark_weights_dark_weights_update_0_write_write_9_stage_95 <= dark_weights_dark_weights_update_0_write_write_9_stage_94;
      dark_weights_dark_weights_update_0_write_write_9_stage_96 <= dark_weights_dark_weights_update_0_write_write_9_stage_95;
      dark_weights_dark_weights_update_0_write_write_9_stage_97 <= dark_weights_dark_weights_update_0_write_write_9_stage_96;
      dark_weights_dark_weights_update_0_write_write_9_stage_98 <= dark_weights_dark_weights_update_0_write_write_9_stage_97;
      dark_weights_dark_weights_update_0_write_write_9_stage_99 <= dark_weights_dark_weights_update_0_write_write_9_stage_98;
      dark_weights_dark_weights_update_0_write_write_9_stage_100 <= dark_weights_dark_weights_update_0_write_write_9_stage_99;
      dark_weights_dark_weights_update_0_write_write_9_stage_101 <= dark_weights_dark_weights_update_0_write_write_9_stage_100;
      dark_weights_dark_weights_update_0_write_write_9_stage_102 <= dark_weights_dark_weights_update_0_write_write_9_stage_101;
      dark_weights_dark_weights_update_0_write_write_9_stage_103 <= dark_weights_dark_weights_update_0_write_write_9_stage_102;
      dark_weights_dark_weights_update_0_write_write_9_stage_104 <= dark_weights_dark_weights_update_0_write_write_9_stage_103;
      dark_weights_dark_weights_update_0_write_write_9_stage_105 <= dark_weights_dark_weights_update_0_write_write_9_stage_104;
      dark_weights_dark_weights_update_0_write_write_9_stage_106 <= dark_weights_dark_weights_update_0_write_write_9_stage_105;
      dark_weights_dark_weights_update_0_write_write_9_stage_107 <= dark_weights_dark_weights_update_0_write_write_9_stage_106;
      dark_weights_dark_weights_update_0_write_write_9_stage_108 <= dark_weights_dark_weights_update_0_write_write_9_stage_107;
      dark_weights_dark_weights_update_0_write_write_9_stage_109 <= dark_weights_dark_weights_update_0_write_write_9_stage_108;
      dark_weights_dark_weights_update_0_write_write_9_stage_110 <= dark_weights_dark_weights_update_0_write_write_9_stage_109;
      dark_weights_dark_weights_update_0_write_write_9_stage_111 <= dark_weights_dark_weights_update_0_write_write_9_stage_110;
      dark_weights_dark_weights_update_0_write_write_9_stage_112 <= dark_weights_dark_weights_update_0_write_write_9_stage_111;
      dark_weights_dark_weights_update_0_write_write_9_stage_113 <= dark_weights_dark_weights_update_0_write_write_9_stage_112;
      dark_weights_dark_weights_update_0_write_write_9_stage_114 <= dark_weights_dark_weights_update_0_write_write_9_stage_113;
      dark_weights_dark_weights_update_0_write_write_9_stage_115 <= dark_weights_dark_weights_update_0_write_write_9_stage_114;
      dark_weights_dark_weights_update_0_write_write_9_stage_116 <= dark_weights_dark_weights_update_0_write_write_9_stage_115;
      dark_weights_dark_weights_update_0_write_write_9_stage_117 <= dark_weights_dark_weights_update_0_write_write_9_stage_116;
      dark_weights_dark_weights_update_0_write_write_9_stage_118 <= dark_weights_dark_weights_update_0_write_write_9_stage_117;
      dark_weights_dark_weights_update_0_write_write_9_stage_119 <= dark_weights_dark_weights_update_0_write_write_9_stage_118;
      dark_weights_dark_weights_update_0_write_write_9_stage_120 <= dark_weights_dark_weights_update_0_write_write_9_stage_119;
      dark_weights_dark_weights_update_0_write_write_9_stage_121 <= dark_weights_dark_weights_update_0_write_write_9_stage_120;
      dark_weights_dark_weights_update_0_write_write_9_stage_122 <= dark_weights_dark_weights_update_0_write_write_9_stage_121;
      dark_weights_dark_weights_update_0_write_write_9_stage_123 <= dark_weights_dark_weights_update_0_write_write_9_stage_122;
      dark_weights_dark_weights_update_0_write_write_9_stage_124 <= dark_weights_dark_weights_update_0_write_write_9_stage_123;
      dark_weights_dark_weights_update_0_write_write_9_stage_125 <= dark_weights_dark_weights_update_0_write_write_9_stage_124;
      dark_weights_dark_weights_update_0_write_write_9_stage_126 <= dark_weights_dark_weights_update_0_write_write_9_stage_125;
      dark_weights_dark_weights_update_0_write_write_9_stage_127 <= dark_weights_dark_weights_update_0_write_write_9_stage_126;
      dark_weights_dark_weights_update_0_write_write_9_stage_128 <= dark_weights_dark_weights_update_0_write_write_9_stage_127;
      dark_weights_dark_weights_update_0_write_write_9_stage_129 <= dark_weights_dark_weights_update_0_write_write_9_stage_128;
      dark_weights_dark_weights_update_0_write_write_9_stage_130 <= dark_weights_dark_weights_update_0_write_write_9_stage_129;
      dark_weights_dark_weights_update_0_write_write_9_stage_131 <= dark_weights_dark_weights_update_0_write_write_9_stage_130;
      dark_weights_dark_weights_update_0_write_write_9_stage_132 <= dark_weights_dark_weights_update_0_write_write_9_stage_131;
      dark_weights_dark_weights_update_0_write_write_9_stage_133 <= dark_weights_dark_weights_update_0_write_write_9_stage_132;
      dark_weights_dark_weights_update_0_write_write_9_stage_134 <= dark_weights_dark_weights_update_0_write_write_9_stage_133;
      dark_weights_dark_weights_update_0_write_write_9_stage_135 <= dark_weights_dark_weights_update_0_write_write_9_stage_134;
      dark_weights_dark_weights_update_0_write_write_9_stage_136 <= dark_weights_dark_weights_update_0_write_write_9_stage_135;
      dark_weights_dark_weights_update_0_write_write_9_stage_137 <= dark_weights_dark_weights_update_0_write_write_9_stage_136;
      dark_weights_dark_weights_update_0_write_write_9_stage_138 <= dark_weights_dark_weights_update_0_write_write_9_stage_137;
      dark_weights_dark_weights_update_0_write_write_9_stage_139 <= dark_weights_dark_weights_update_0_write_write_9_stage_138;
      dark_weights_dark_weights_update_0_write_write_9_stage_140 <= dark_weights_dark_weights_update_0_write_write_9_stage_139;
      dark_weights_dark_weights_update_0_write_write_9_stage_141 <= dark_weights_dark_weights_update_0_write_write_9_stage_140;
      dark_weights_dark_weights_update_0_write_write_9_stage_142 <= dark_weights_dark_weights_update_0_write_write_9_stage_141;
      dark_weights_dark_weights_update_0_write_write_9_stage_143 <= dark_weights_dark_weights_update_0_write_write_9_stage_142;
      dark_weights_dark_weights_update_0_write_write_9_stage_144 <= dark_weights_dark_weights_update_0_write_write_9_stage_143;
      dark_weights_dark_weights_update_0_write_write_9_stage_145 <= dark_weights_dark_weights_update_0_write_write_9_stage_144;
      dark_weights_dark_weights_update_0_write_write_9_stage_146 <= dark_weights_dark_weights_update_0_write_write_9_stage_145;
      dark_weights_dark_weights_update_0_write_write_9_stage_147 <= dark_weights_dark_weights_update_0_write_write_9_stage_146;
      dark_weights_dark_weights_update_0_write_write_9_stage_148 <= dark_weights_dark_weights_update_0_write_write_9_stage_147;
      dark_weights_dark_weights_update_0_write_write_9_stage_149 <= dark_weights_dark_weights_update_0_write_write_9_stage_148;
      dark_weights_dark_weights_update_0_write_write_9_stage_150 <= dark_weights_dark_weights_update_0_write_write_9_stage_149;
      dark_weights_dark_weights_update_0_write_write_9_stage_151 <= dark_weights_dark_weights_update_0_write_write_9_stage_150;
      dark_weights_dark_weights_update_0_write_write_9_stage_152 <= dark_weights_dark_weights_update_0_write_write_9_stage_151;
      dark_weights_dark_weights_update_0_write_write_9_stage_153 <= dark_weights_dark_weights_update_0_write_write_9_stage_152;
      dark_weights_dark_weights_update_0_write_write_9_stage_154 <= dark_weights_dark_weights_update_0_write_write_9_stage_153;
      dark_weights_dark_weights_update_0_write_write_9_stage_155 <= dark_weights_dark_weights_update_0_write_write_9_stage_154;
      dark_weights_dark_weights_update_0_write_write_9_stage_156 <= dark_weights_dark_weights_update_0_write_write_9_stage_155;
      dark_weights_dark_weights_update_0_write_write_9_stage_157 <= dark_weights_dark_weights_update_0_write_write_9_stage_156;
      dark_weights_dark_weights_update_0_write_write_9_stage_158 <= dark_weights_dark_weights_update_0_write_write_9_stage_157;
      dark_weights_dark_weights_update_0_write_write_9_stage_159 <= dark_weights_dark_weights_update_0_write_write_9_stage_158;
      dark_weights_dark_weights_update_0_write_write_9_stage_160 <= dark_weights_dark_weights_update_0_write_write_9_stage_159;
      dark_weights_dark_weights_update_0_write_write_9_stage_161 <= dark_weights_dark_weights_update_0_write_write_9_stage_160;
      dark_weights_dark_weights_update_0_write_write_9_stage_162 <= dark_weights_dark_weights_update_0_write_write_9_stage_161;
      dark_weights_dark_weights_update_0_write_write_9_stage_163 <= dark_weights_dark_weights_update_0_write_write_9_stage_162;
      dark_weights_dark_weights_update_0_write_write_9_stage_164 <= dark_weights_dark_weights_update_0_write_write_9_stage_163;
      dark_weights_dark_weights_update_0_write_write_9_stage_165 <= dark_weights_dark_weights_update_0_write_write_9_stage_164;
      dark_weights_dark_weights_update_0_write_write_9_stage_166 <= dark_weights_dark_weights_update_0_write_write_9_stage_165;
      dark_weights_dark_weights_update_0_write_write_9_stage_167 <= dark_weights_dark_weights_update_0_write_write_9_stage_166;
      dark_weights_dark_weights_update_0_write_write_9_stage_168 <= dark_weights_dark_weights_update_0_write_write_9_stage_167;
      dark_weights_dark_weights_update_0_write_write_9_stage_169 <= dark_weights_dark_weights_update_0_write_write_9_stage_168;
      dark_weights_dark_weights_update_0_write_write_9_stage_170 <= dark_weights_dark_weights_update_0_write_write_9_stage_169;
      dark_weights_dark_weights_update_0_write_write_9_stage_171 <= dark_weights_dark_weights_update_0_write_write_9_stage_170;
      dark_weights_dark_weights_update_0_write_write_9_stage_172 <= dark_weights_dark_weights_update_0_write_write_9_stage_171;
      dark_weights_dark_weights_update_0_write_write_9_stage_173 <= dark_weights_dark_weights_update_0_write_write_9_stage_172;
      dark_weights_dark_weights_update_0_write_write_9_stage_174 <= dark_weights_dark_weights_update_0_write_write_9_stage_173;
      dark_weights_dark_weights_update_0_write_write_9_stage_175 <= dark_weights_dark_weights_update_0_write_write_9_stage_174;
      dark_weights_dark_weights_update_0_write_write_9_stage_176 <= dark_weights_dark_weights_update_0_write_write_9_stage_175;
      dark_weights_dark_weights_update_0_write_write_9_stage_177 <= dark_weights_dark_weights_update_0_write_write_9_stage_176;
      dark_weights_dark_weights_update_0_write_write_9_stage_178 <= dark_weights_dark_weights_update_0_write_write_9_stage_177;
      dark_weights_dark_weights_update_0_write_write_9_stage_179 <= dark_weights_dark_weights_update_0_write_write_9_stage_178;
      dark_weights_dark_weights_update_0_write_write_9_stage_180 <= dark_weights_dark_weights_update_0_write_write_9_stage_179;
      dark_weights_dark_weights_update_0_write_write_9_stage_181 <= dark_weights_dark_weights_update_0_write_write_9_stage_180;
      dark_weights_normed_gauss_blur_2_update_0_stage_86 <= dark_weights_normed_gauss_blur_2_update_0;
      dark_weights_normed_gauss_blur_2_update_0_stage_87 <= dark_weights_normed_gauss_blur_2_update_0_stage_86;
      dark_weights_normed_gauss_blur_2_update_0_stage_88 <= dark_weights_normed_gauss_blur_2_update_0_stage_87;
      dark_weights_normed_gauss_blur_2_update_0_stage_89 <= dark_weights_normed_gauss_blur_2_update_0_stage_88;
      dark_weights_normed_gauss_blur_2_update_0_stage_90 <= dark_weights_normed_gauss_blur_2_update_0_stage_89;
      dark_weights_normed_gauss_blur_2_update_0_stage_91 <= dark_weights_normed_gauss_blur_2_update_0_stage_90;
      dark_weights_normed_gauss_blur_2_update_0_stage_92 <= dark_weights_normed_gauss_blur_2_update_0_stage_91;
      dark_weights_normed_gauss_blur_2_update_0_stage_93 <= dark_weights_normed_gauss_blur_2_update_0_stage_92;
      dark_weights_normed_gauss_blur_2_update_0_stage_94 <= dark_weights_normed_gauss_blur_2_update_0_stage_93;
      dark_weights_normed_gauss_blur_2_update_0_stage_95 <= dark_weights_normed_gauss_blur_2_update_0_stage_94;
      dark_weights_normed_gauss_blur_2_update_0_stage_96 <= dark_weights_normed_gauss_blur_2_update_0_stage_95;
      dark_weights_normed_gauss_blur_2_update_0_stage_97 <= dark_weights_normed_gauss_blur_2_update_0_stage_96;
      dark_weights_normed_gauss_blur_2_update_0_stage_98 <= dark_weights_normed_gauss_blur_2_update_0_stage_97;
      dark_weights_normed_gauss_blur_2_update_0_stage_99 <= dark_weights_normed_gauss_blur_2_update_0_stage_98;
      dark_weights_normed_gauss_blur_2_update_0_stage_100 <= dark_weights_normed_gauss_blur_2_update_0_stage_99;
      dark_weights_normed_gauss_blur_2_update_0_stage_101 <= dark_weights_normed_gauss_blur_2_update_0_stage_100;
      dark_weights_normed_gauss_blur_2_update_0_stage_102 <= dark_weights_normed_gauss_blur_2_update_0_stage_101;
      dark_weights_normed_gauss_blur_2_update_0_stage_103 <= dark_weights_normed_gauss_blur_2_update_0_stage_102;
      dark_weights_normed_gauss_blur_2_update_0_stage_104 <= dark_weights_normed_gauss_blur_2_update_0_stage_103;
      dark_weights_normed_gauss_blur_2_update_0_stage_105 <= dark_weights_normed_gauss_blur_2_update_0_stage_104;
      dark_weights_normed_gauss_blur_2_update_0_stage_106 <= dark_weights_normed_gauss_blur_2_update_0_stage_105;
      dark_weights_normed_gauss_blur_2_update_0_stage_107 <= dark_weights_normed_gauss_blur_2_update_0_stage_106;
      dark_weights_normed_gauss_blur_2_update_0_stage_108 <= dark_weights_normed_gauss_blur_2_update_0_stage_107;
      dark_weights_normed_gauss_blur_2_update_0_stage_109 <= dark_weights_normed_gauss_blur_2_update_0_stage_108;
      dark_weights_normed_gauss_blur_2_update_0_stage_110 <= dark_weights_normed_gauss_blur_2_update_0_stage_109;
      dark_weights_normed_gauss_blur_2_update_0_stage_111 <= dark_weights_normed_gauss_blur_2_update_0_stage_110;
      dark_weights_normed_gauss_blur_2_update_0_stage_112 <= dark_weights_normed_gauss_blur_2_update_0_stage_111;
      dark_weights_normed_gauss_blur_2_update_0_stage_113 <= dark_weights_normed_gauss_blur_2_update_0_stage_112;
      dark_weights_normed_gauss_blur_2_update_0_stage_114 <= dark_weights_normed_gauss_blur_2_update_0_stage_113;
      dark_weights_normed_gauss_blur_2_update_0_stage_115 <= dark_weights_normed_gauss_blur_2_update_0_stage_114;
      dark_weights_normed_gauss_blur_2_update_0_stage_116 <= dark_weights_normed_gauss_blur_2_update_0_stage_115;
      dark_weights_normed_gauss_blur_2_update_0_stage_117 <= dark_weights_normed_gauss_blur_2_update_0_stage_116;
      dark_weights_normed_gauss_blur_2_update_0_stage_118 <= dark_weights_normed_gauss_blur_2_update_0_stage_117;
      dark_weights_normed_gauss_blur_2_update_0_stage_119 <= dark_weights_normed_gauss_blur_2_update_0_stage_118;
      dark_weights_normed_gauss_blur_2_update_0_stage_120 <= dark_weights_normed_gauss_blur_2_update_0_stage_119;
      dark_weights_normed_gauss_blur_2_update_0_stage_121 <= dark_weights_normed_gauss_blur_2_update_0_stage_120;
      dark_weights_normed_gauss_blur_2_update_0_stage_122 <= dark_weights_normed_gauss_blur_2_update_0_stage_121;
      dark_weights_normed_gauss_blur_2_update_0_stage_123 <= dark_weights_normed_gauss_blur_2_update_0_stage_122;
      dark_weights_normed_gauss_blur_2_update_0_stage_124 <= dark_weights_normed_gauss_blur_2_update_0_stage_123;
      dark_weights_normed_gauss_blur_2_update_0_stage_125 <= dark_weights_normed_gauss_blur_2_update_0_stage_124;
      dark_weights_normed_gauss_blur_2_update_0_stage_126 <= dark_weights_normed_gauss_blur_2_update_0_stage_125;
      dark_weights_normed_gauss_blur_2_update_0_stage_127 <= dark_weights_normed_gauss_blur_2_update_0_stage_126;
      dark_weights_normed_gauss_blur_2_update_0_stage_128 <= dark_weights_normed_gauss_blur_2_update_0_stage_127;
      dark_weights_normed_gauss_blur_2_update_0_stage_129 <= dark_weights_normed_gauss_blur_2_update_0_stage_128;
      dark_weights_normed_gauss_blur_2_update_0_stage_130 <= dark_weights_normed_gauss_blur_2_update_0_stage_129;
      dark_weights_normed_gauss_blur_2_update_0_stage_131 <= dark_weights_normed_gauss_blur_2_update_0_stage_130;
      dark_weights_normed_gauss_blur_2_update_0_stage_132 <= dark_weights_normed_gauss_blur_2_update_0_stage_131;
      dark_weights_normed_gauss_blur_2_update_0_stage_133 <= dark_weights_normed_gauss_blur_2_update_0_stage_132;
      dark_weights_normed_gauss_blur_2_update_0_stage_134 <= dark_weights_normed_gauss_blur_2_update_0_stage_133;
      dark_weights_normed_gauss_blur_2_update_0_stage_135 <= dark_weights_normed_gauss_blur_2_update_0_stage_134;
      dark_weights_normed_gauss_blur_2_update_0_stage_136 <= dark_weights_normed_gauss_blur_2_update_0_stage_135;
      dark_weights_normed_gauss_blur_2_update_0_stage_137 <= dark_weights_normed_gauss_blur_2_update_0_stage_136;
      dark_weights_normed_gauss_blur_2_update_0_stage_138 <= dark_weights_normed_gauss_blur_2_update_0_stage_137;
      dark_weights_normed_gauss_blur_2_update_0_stage_139 <= dark_weights_normed_gauss_blur_2_update_0_stage_138;
      dark_weights_normed_gauss_blur_2_update_0_stage_140 <= dark_weights_normed_gauss_blur_2_update_0_stage_139;
      dark_weights_normed_gauss_blur_2_update_0_stage_141 <= dark_weights_normed_gauss_blur_2_update_0_stage_140;
      dark_weights_normed_gauss_blur_2_update_0_stage_142 <= dark_weights_normed_gauss_blur_2_update_0_stage_141;
      dark_weights_normed_gauss_blur_2_update_0_stage_143 <= dark_weights_normed_gauss_blur_2_update_0_stage_142;
      dark_weights_normed_gauss_blur_2_update_0_stage_144 <= dark_weights_normed_gauss_blur_2_update_0_stage_143;
      dark_weights_normed_gauss_blur_2_update_0_stage_145 <= dark_weights_normed_gauss_blur_2_update_0_stage_144;
      dark_weights_normed_gauss_blur_2_update_0_stage_146 <= dark_weights_normed_gauss_blur_2_update_0_stage_145;
      dark_weights_normed_gauss_blur_2_update_0_stage_147 <= dark_weights_normed_gauss_blur_2_update_0_stage_146;
      dark_weights_normed_gauss_blur_2_update_0_stage_148 <= dark_weights_normed_gauss_blur_2_update_0_stage_147;
      dark_weights_normed_gauss_blur_2_update_0_stage_149 <= dark_weights_normed_gauss_blur_2_update_0_stage_148;
      dark_weights_normed_gauss_blur_2_update_0_stage_150 <= dark_weights_normed_gauss_blur_2_update_0_stage_149;
      dark_weights_normed_gauss_blur_2_update_0_stage_151 <= dark_weights_normed_gauss_blur_2_update_0_stage_150;
      dark_weights_normed_gauss_blur_2_update_0_stage_152 <= dark_weights_normed_gauss_blur_2_update_0_stage_151;
      dark_weights_normed_gauss_blur_2_update_0_stage_153 <= dark_weights_normed_gauss_blur_2_update_0_stage_152;
      dark_weights_normed_gauss_blur_2_update_0_stage_154 <= dark_weights_normed_gauss_blur_2_update_0_stage_153;
      dark_weights_normed_gauss_blur_2_update_0_stage_155 <= dark_weights_normed_gauss_blur_2_update_0_stage_154;
      dark_weights_normed_gauss_blur_2_update_0_stage_156 <= dark_weights_normed_gauss_blur_2_update_0_stage_155;
      dark_weights_normed_gauss_blur_2_update_0_stage_157 <= dark_weights_normed_gauss_blur_2_update_0_stage_156;
      dark_weights_normed_gauss_blur_2_update_0_stage_158 <= dark_weights_normed_gauss_blur_2_update_0_stage_157;
      dark_weights_normed_gauss_blur_2_update_0_stage_159 <= dark_weights_normed_gauss_blur_2_update_0_stage_158;
      dark_weights_normed_gauss_blur_2_update_0_stage_160 <= dark_weights_normed_gauss_blur_2_update_0_stage_159;
      dark_weights_normed_gauss_blur_2_update_0_stage_161 <= dark_weights_normed_gauss_blur_2_update_0_stage_160;
      dark_weights_normed_gauss_blur_2_update_0_stage_162 <= dark_weights_normed_gauss_blur_2_update_0_stage_161;
      dark_weights_normed_gauss_blur_2_update_0_stage_163 <= dark_weights_normed_gauss_blur_2_update_0_stage_162;
      dark_weights_normed_gauss_blur_2_update_0_stage_164 <= dark_weights_normed_gauss_blur_2_update_0_stage_163;
      dark_weights_normed_gauss_blur_2_update_0_stage_165 <= dark_weights_normed_gauss_blur_2_update_0_stage_164;
      dark_weights_normed_gauss_blur_2_update_0_stage_166 <= dark_weights_normed_gauss_blur_2_update_0_stage_165;
      dark_weights_normed_gauss_blur_2_update_0_stage_167 <= dark_weights_normed_gauss_blur_2_update_0_stage_166;
      dark_weights_normed_gauss_blur_2_update_0_stage_168 <= dark_weights_normed_gauss_blur_2_update_0_stage_167;
      dark_weights_normed_gauss_blur_2_update_0_stage_169 <= dark_weights_normed_gauss_blur_2_update_0_stage_168;
      dark_weights_normed_gauss_blur_2_update_0_stage_170 <= dark_weights_normed_gauss_blur_2_update_0_stage_169;
      dark_weights_normed_gauss_blur_2_update_0_stage_171 <= dark_weights_normed_gauss_blur_2_update_0_stage_170;
      dark_weights_normed_gauss_blur_2_update_0_stage_172 <= dark_weights_normed_gauss_blur_2_update_0_stage_171;
      dark_weights_normed_gauss_blur_2_update_0_stage_173 <= dark_weights_normed_gauss_blur_2_update_0_stage_172;
      dark_weights_normed_gauss_blur_2_update_0_stage_174 <= dark_weights_normed_gauss_blur_2_update_0_stage_173;
      dark_weights_normed_gauss_blur_2_update_0_stage_175 <= dark_weights_normed_gauss_blur_2_update_0_stage_174;
      dark_weights_normed_gauss_blur_2_update_0_stage_176 <= dark_weights_normed_gauss_blur_2_update_0_stage_175;
      dark_weights_normed_gauss_blur_2_update_0_stage_177 <= dark_weights_normed_gauss_blur_2_update_0_stage_176;
      dark_weights_normed_gauss_blur_2_update_0_stage_178 <= dark_weights_normed_gauss_blur_2_update_0_stage_177;
      dark_weights_normed_gauss_blur_2_update_0_stage_179 <= dark_weights_normed_gauss_blur_2_update_0_stage_178;
      dark_weights_normed_gauss_blur_2_update_0_stage_180 <= dark_weights_normed_gauss_blur_2_update_0_stage_179;
      dark_weights_normed_gauss_blur_2_update_0_stage_181 <= dark_weights_normed_gauss_blur_2_update_0_stage_180;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_171 <= final_merged_2_final_merged_1_update_0_read_read_120;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_172 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_171;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_173 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_172;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_174 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_173;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_175 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_174;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_176 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_175;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_177 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_176;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_178 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_177;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_179 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_178;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_180 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_179;
      final_merged_2_final_merged_1_update_0_read_read_120_stage_181 <= final_merged_2_final_merged_1_update_0_read_read_120_stage_180;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_87 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_88 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_87;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_89 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_88;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_90 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_89;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_91 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_90;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_92 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_91;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_93 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_92;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_94 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_93;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_95 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_94;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_96 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_95;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_97 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_96;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_98 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_97;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_99 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_98;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_100 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_99;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_101 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_100;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_102 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_101;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_103 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_102;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_104 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_103;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_105 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_104;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_106 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_105;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_107 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_106;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_108 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_107;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_109 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_108;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_110 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_109;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_111 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_110;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_112 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_111;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_113 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_112;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_114 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_113;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_115 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_114;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_116 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_115;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_117 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_116;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_118 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_117;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_119 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_118;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_120 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_119;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_121 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_120;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_122 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_121;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_123 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_122;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_124 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_123;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_125 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_124;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_126 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_125;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_127 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_126;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_128 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_127;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_129 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_128;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_130 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_129;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_131 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_130;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_132 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_131;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_133 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_132;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_134 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_133;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_135 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_134;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_136 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_135;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_137 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_136;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_138 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_137;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_139 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_138;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_140 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_139;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_141 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_140;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_142 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_141;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_143 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_142;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_144 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_143;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_145 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_144;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_146 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_145;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_147 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_146;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_148 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_147;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_149 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_148;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_150 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_149;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_151 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_150;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_152 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_151;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_153 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_152;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_154 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_153;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_155 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_154;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_156 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_155;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_157 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_156;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_158 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_157;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_159 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_158;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_160 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_159;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_161 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_160;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_162 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_161;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_163 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_162;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_164 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_163;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_165 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_164;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_166 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_165;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_167 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_166;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_168 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_167;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_169 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_168;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_170 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_169;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_171 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_170;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_172 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_171;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_173 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_172;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_174 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_173;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_175 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_174;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_176 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_175;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_177 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_176;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_178 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_177;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_179 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_178;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_180 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_179;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_181 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58_stage_180;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_172 <= fused_level_1_final_merged_1_update_0_read_read_121;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_173 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_172;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_174 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_173;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_175 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_174;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_176 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_175;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_177 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_176;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_178 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_177;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_179 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_178;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_180 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_179;
      fused_level_1_final_merged_1_update_0_read_read_121_stage_181 <= fused_level_1_final_merged_1_update_0_read_read_121_stage_180;
      final_merged_1_update_0_stage_173 <= final_merged_1_update_0;
      final_merged_1_update_0_stage_174 <= final_merged_1_update_0_stage_173;
      final_merged_1_update_0_stage_175 <= final_merged_1_update_0_stage_174;
      final_merged_1_update_0_stage_176 <= final_merged_1_update_0_stage_175;
      final_merged_1_update_0_stage_177 <= final_merged_1_update_0_stage_176;
      final_merged_1_update_0_stage_178 <= final_merged_1_update_0_stage_177;
      final_merged_1_update_0_stage_179 <= final_merged_1_update_0_stage_178;
      final_merged_1_update_0_stage_180 <= final_merged_1_update_0_stage_179;
      final_merged_1_update_0_stage_181 <= final_merged_1_update_0_stage_180;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_174 <= final_merged_1_final_merged_1_update_0_write_write_122;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_175 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_174;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_176 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_175;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_177 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_176;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_178 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_177;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_179 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_178;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_180 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_179;
      final_merged_1_final_merged_1_update_0_write_write_122_stage_181 <= final_merged_1_final_merged_1_update_0_write_write_122_stage_180;
      in_in_update_0_write_write_1_stage_4 <= in_in_update_0_write_write_1;
      in_in_update_0_write_write_1_stage_5 <= in_in_update_0_write_write_1_stage_4;
      in_in_update_0_write_write_1_stage_6 <= in_in_update_0_write_write_1_stage_5;
      in_in_update_0_write_write_1_stage_7 <= in_in_update_0_write_write_1_stage_6;
      in_in_update_0_write_write_1_stage_8 <= in_in_update_0_write_write_1_stage_7;
      in_in_update_0_write_write_1_stage_9 <= in_in_update_0_write_write_1_stage_8;
      in_in_update_0_write_write_1_stage_10 <= in_in_update_0_write_write_1_stage_9;
      in_in_update_0_write_write_1_stage_11 <= in_in_update_0_write_write_1_stage_10;
      in_in_update_0_write_write_1_stage_12 <= in_in_update_0_write_write_1_stage_11;
      in_in_update_0_write_write_1_stage_13 <= in_in_update_0_write_write_1_stage_12;
      in_in_update_0_write_write_1_stage_14 <= in_in_update_0_write_write_1_stage_13;
      in_in_update_0_write_write_1_stage_15 <= in_in_update_0_write_write_1_stage_14;
      in_in_update_0_write_write_1_stage_16 <= in_in_update_0_write_write_1_stage_15;
      in_in_update_0_write_write_1_stage_17 <= in_in_update_0_write_write_1_stage_16;
      in_in_update_0_write_write_1_stage_18 <= in_in_update_0_write_write_1_stage_17;
      in_in_update_0_write_write_1_stage_19 <= in_in_update_0_write_write_1_stage_18;
      in_in_update_0_write_write_1_stage_20 <= in_in_update_0_write_write_1_stage_19;
      in_in_update_0_write_write_1_stage_21 <= in_in_update_0_write_write_1_stage_20;
      in_in_update_0_write_write_1_stage_22 <= in_in_update_0_write_write_1_stage_21;
      in_in_update_0_write_write_1_stage_23 <= in_in_update_0_write_write_1_stage_22;
      in_in_update_0_write_write_1_stage_24 <= in_in_update_0_write_write_1_stage_23;
      in_in_update_0_write_write_1_stage_25 <= in_in_update_0_write_write_1_stage_24;
      in_in_update_0_write_write_1_stage_26 <= in_in_update_0_write_write_1_stage_25;
      in_in_update_0_write_write_1_stage_27 <= in_in_update_0_write_write_1_stage_26;
      in_in_update_0_write_write_1_stage_28 <= in_in_update_0_write_write_1_stage_27;
      in_in_update_0_write_write_1_stage_29 <= in_in_update_0_write_write_1_stage_28;
      in_in_update_0_write_write_1_stage_30 <= in_in_update_0_write_write_1_stage_29;
      in_in_update_0_write_write_1_stage_31 <= in_in_update_0_write_write_1_stage_30;
      in_in_update_0_write_write_1_stage_32 <= in_in_update_0_write_write_1_stage_31;
      in_in_update_0_write_write_1_stage_33 <= in_in_update_0_write_write_1_stage_32;
      in_in_update_0_write_write_1_stage_34 <= in_in_update_0_write_write_1_stage_33;
      in_in_update_0_write_write_1_stage_35 <= in_in_update_0_write_write_1_stage_34;
      in_in_update_0_write_write_1_stage_36 <= in_in_update_0_write_write_1_stage_35;
      in_in_update_0_write_write_1_stage_37 <= in_in_update_0_write_write_1_stage_36;
      in_in_update_0_write_write_1_stage_38 <= in_in_update_0_write_write_1_stage_37;
      in_in_update_0_write_write_1_stage_39 <= in_in_update_0_write_write_1_stage_38;
      in_in_update_0_write_write_1_stage_40 <= in_in_update_0_write_write_1_stage_39;
      in_in_update_0_write_write_1_stage_41 <= in_in_update_0_write_write_1_stage_40;
      in_in_update_0_write_write_1_stage_42 <= in_in_update_0_write_write_1_stage_41;
      in_in_update_0_write_write_1_stage_43 <= in_in_update_0_write_write_1_stage_42;
      in_in_update_0_write_write_1_stage_44 <= in_in_update_0_write_write_1_stage_43;
      in_in_update_0_write_write_1_stage_45 <= in_in_update_0_write_write_1_stage_44;
      in_in_update_0_write_write_1_stage_46 <= in_in_update_0_write_write_1_stage_45;
      in_in_update_0_write_write_1_stage_47 <= in_in_update_0_write_write_1_stage_46;
      in_in_update_0_write_write_1_stage_48 <= in_in_update_0_write_write_1_stage_47;
      in_in_update_0_write_write_1_stage_49 <= in_in_update_0_write_write_1_stage_48;
      in_in_update_0_write_write_1_stage_50 <= in_in_update_0_write_write_1_stage_49;
      in_in_update_0_write_write_1_stage_51 <= in_in_update_0_write_write_1_stage_50;
      in_in_update_0_write_write_1_stage_52 <= in_in_update_0_write_write_1_stage_51;
      in_in_update_0_write_write_1_stage_53 <= in_in_update_0_write_write_1_stage_52;
      in_in_update_0_write_write_1_stage_54 <= in_in_update_0_write_write_1_stage_53;
      in_in_update_0_write_write_1_stage_55 <= in_in_update_0_write_write_1_stage_54;
      in_in_update_0_write_write_1_stage_56 <= in_in_update_0_write_write_1_stage_55;
      in_in_update_0_write_write_1_stage_57 <= in_in_update_0_write_write_1_stage_56;
      in_in_update_0_write_write_1_stage_58 <= in_in_update_0_write_write_1_stage_57;
      in_in_update_0_write_write_1_stage_59 <= in_in_update_0_write_write_1_stage_58;
      in_in_update_0_write_write_1_stage_60 <= in_in_update_0_write_write_1_stage_59;
      in_in_update_0_write_write_1_stage_61 <= in_in_update_0_write_write_1_stage_60;
      in_in_update_0_write_write_1_stage_62 <= in_in_update_0_write_write_1_stage_61;
      in_in_update_0_write_write_1_stage_63 <= in_in_update_0_write_write_1_stage_62;
      in_in_update_0_write_write_1_stage_64 <= in_in_update_0_write_write_1_stage_63;
      in_in_update_0_write_write_1_stage_65 <= in_in_update_0_write_write_1_stage_64;
      in_in_update_0_write_write_1_stage_66 <= in_in_update_0_write_write_1_stage_65;
      in_in_update_0_write_write_1_stage_67 <= in_in_update_0_write_write_1_stage_66;
      in_in_update_0_write_write_1_stage_68 <= in_in_update_0_write_write_1_stage_67;
      in_in_update_0_write_write_1_stage_69 <= in_in_update_0_write_write_1_stage_68;
      in_in_update_0_write_write_1_stage_70 <= in_in_update_0_write_write_1_stage_69;
      in_in_update_0_write_write_1_stage_71 <= in_in_update_0_write_write_1_stage_70;
      in_in_update_0_write_write_1_stage_72 <= in_in_update_0_write_write_1_stage_71;
      in_in_update_0_write_write_1_stage_73 <= in_in_update_0_write_write_1_stage_72;
      in_in_update_0_write_write_1_stage_74 <= in_in_update_0_write_write_1_stage_73;
      in_in_update_0_write_write_1_stage_75 <= in_in_update_0_write_write_1_stage_74;
      in_in_update_0_write_write_1_stage_76 <= in_in_update_0_write_write_1_stage_75;
      in_in_update_0_write_write_1_stage_77 <= in_in_update_0_write_write_1_stage_76;
      in_in_update_0_write_write_1_stage_78 <= in_in_update_0_write_write_1_stage_77;
      in_in_update_0_write_write_1_stage_79 <= in_in_update_0_write_write_1_stage_78;
      in_in_update_0_write_write_1_stage_80 <= in_in_update_0_write_write_1_stage_79;
      in_in_update_0_write_write_1_stage_81 <= in_in_update_0_write_write_1_stage_80;
      in_in_update_0_write_write_1_stage_82 <= in_in_update_0_write_write_1_stage_81;
      in_in_update_0_write_write_1_stage_83 <= in_in_update_0_write_write_1_stage_82;
      in_in_update_0_write_write_1_stage_84 <= in_in_update_0_write_write_1_stage_83;
      in_in_update_0_write_write_1_stage_85 <= in_in_update_0_write_write_1_stage_84;
      in_in_update_0_write_write_1_stage_86 <= in_in_update_0_write_write_1_stage_85;
      in_in_update_0_write_write_1_stage_87 <= in_in_update_0_write_write_1_stage_86;
      in_in_update_0_write_write_1_stage_88 <= in_in_update_0_write_write_1_stage_87;
      in_in_update_0_write_write_1_stage_89 <= in_in_update_0_write_write_1_stage_88;
      in_in_update_0_write_write_1_stage_90 <= in_in_update_0_write_write_1_stage_89;
      in_in_update_0_write_write_1_stage_91 <= in_in_update_0_write_write_1_stage_90;
      in_in_update_0_write_write_1_stage_92 <= in_in_update_0_write_write_1_stage_91;
      in_in_update_0_write_write_1_stage_93 <= in_in_update_0_write_write_1_stage_92;
      in_in_update_0_write_write_1_stage_94 <= in_in_update_0_write_write_1_stage_93;
      in_in_update_0_write_write_1_stage_95 <= in_in_update_0_write_write_1_stage_94;
      in_in_update_0_write_write_1_stage_96 <= in_in_update_0_write_write_1_stage_95;
      in_in_update_0_write_write_1_stage_97 <= in_in_update_0_write_write_1_stage_96;
      in_in_update_0_write_write_1_stage_98 <= in_in_update_0_write_write_1_stage_97;
      in_in_update_0_write_write_1_stage_99 <= in_in_update_0_write_write_1_stage_98;
      in_in_update_0_write_write_1_stage_100 <= in_in_update_0_write_write_1_stage_99;
      in_in_update_0_write_write_1_stage_101 <= in_in_update_0_write_write_1_stage_100;
      in_in_update_0_write_write_1_stage_102 <= in_in_update_0_write_write_1_stage_101;
      in_in_update_0_write_write_1_stage_103 <= in_in_update_0_write_write_1_stage_102;
      in_in_update_0_write_write_1_stage_104 <= in_in_update_0_write_write_1_stage_103;
      in_in_update_0_write_write_1_stage_105 <= in_in_update_0_write_write_1_stage_104;
      in_in_update_0_write_write_1_stage_106 <= in_in_update_0_write_write_1_stage_105;
      in_in_update_0_write_write_1_stage_107 <= in_in_update_0_write_write_1_stage_106;
      in_in_update_0_write_write_1_stage_108 <= in_in_update_0_write_write_1_stage_107;
      in_in_update_0_write_write_1_stage_109 <= in_in_update_0_write_write_1_stage_108;
      in_in_update_0_write_write_1_stage_110 <= in_in_update_0_write_write_1_stage_109;
      in_in_update_0_write_write_1_stage_111 <= in_in_update_0_write_write_1_stage_110;
      in_in_update_0_write_write_1_stage_112 <= in_in_update_0_write_write_1_stage_111;
      in_in_update_0_write_write_1_stage_113 <= in_in_update_0_write_write_1_stage_112;
      in_in_update_0_write_write_1_stage_114 <= in_in_update_0_write_write_1_stage_113;
      in_in_update_0_write_write_1_stage_115 <= in_in_update_0_write_write_1_stage_114;
      in_in_update_0_write_write_1_stage_116 <= in_in_update_0_write_write_1_stage_115;
      in_in_update_0_write_write_1_stage_117 <= in_in_update_0_write_write_1_stage_116;
      in_in_update_0_write_write_1_stage_118 <= in_in_update_0_write_write_1_stage_117;
      in_in_update_0_write_write_1_stage_119 <= in_in_update_0_write_write_1_stage_118;
      in_in_update_0_write_write_1_stage_120 <= in_in_update_0_write_write_1_stage_119;
      in_in_update_0_write_write_1_stage_121 <= in_in_update_0_write_write_1_stage_120;
      in_in_update_0_write_write_1_stage_122 <= in_in_update_0_write_write_1_stage_121;
      in_in_update_0_write_write_1_stage_123 <= in_in_update_0_write_write_1_stage_122;
      in_in_update_0_write_write_1_stage_124 <= in_in_update_0_write_write_1_stage_123;
      in_in_update_0_write_write_1_stage_125 <= in_in_update_0_write_write_1_stage_124;
      in_in_update_0_write_write_1_stage_126 <= in_in_update_0_write_write_1_stage_125;
      in_in_update_0_write_write_1_stage_127 <= in_in_update_0_write_write_1_stage_126;
      in_in_update_0_write_write_1_stage_128 <= in_in_update_0_write_write_1_stage_127;
      in_in_update_0_write_write_1_stage_129 <= in_in_update_0_write_write_1_stage_128;
      in_in_update_0_write_write_1_stage_130 <= in_in_update_0_write_write_1_stage_129;
      in_in_update_0_write_write_1_stage_131 <= in_in_update_0_write_write_1_stage_130;
      in_in_update_0_write_write_1_stage_132 <= in_in_update_0_write_write_1_stage_131;
      in_in_update_0_write_write_1_stage_133 <= in_in_update_0_write_write_1_stage_132;
      in_in_update_0_write_write_1_stage_134 <= in_in_update_0_write_write_1_stage_133;
      in_in_update_0_write_write_1_stage_135 <= in_in_update_0_write_write_1_stage_134;
      in_in_update_0_write_write_1_stage_136 <= in_in_update_0_write_write_1_stage_135;
      in_in_update_0_write_write_1_stage_137 <= in_in_update_0_write_write_1_stage_136;
      in_in_update_0_write_write_1_stage_138 <= in_in_update_0_write_write_1_stage_137;
      in_in_update_0_write_write_1_stage_139 <= in_in_update_0_write_write_1_stage_138;
      in_in_update_0_write_write_1_stage_140 <= in_in_update_0_write_write_1_stage_139;
      in_in_update_0_write_write_1_stage_141 <= in_in_update_0_write_write_1_stage_140;
      in_in_update_0_write_write_1_stage_142 <= in_in_update_0_write_write_1_stage_141;
      in_in_update_0_write_write_1_stage_143 <= in_in_update_0_write_write_1_stage_142;
      in_in_update_0_write_write_1_stage_144 <= in_in_update_0_write_write_1_stage_143;
      in_in_update_0_write_write_1_stage_145 <= in_in_update_0_write_write_1_stage_144;
      in_in_update_0_write_write_1_stage_146 <= in_in_update_0_write_write_1_stage_145;
      in_in_update_0_write_write_1_stage_147 <= in_in_update_0_write_write_1_stage_146;
      in_in_update_0_write_write_1_stage_148 <= in_in_update_0_write_write_1_stage_147;
      in_in_update_0_write_write_1_stage_149 <= in_in_update_0_write_write_1_stage_148;
      in_in_update_0_write_write_1_stage_150 <= in_in_update_0_write_write_1_stage_149;
      in_in_update_0_write_write_1_stage_151 <= in_in_update_0_write_write_1_stage_150;
      in_in_update_0_write_write_1_stage_152 <= in_in_update_0_write_write_1_stage_151;
      in_in_update_0_write_write_1_stage_153 <= in_in_update_0_write_write_1_stage_152;
      in_in_update_0_write_write_1_stage_154 <= in_in_update_0_write_write_1_stage_153;
      in_in_update_0_write_write_1_stage_155 <= in_in_update_0_write_write_1_stage_154;
      in_in_update_0_write_write_1_stage_156 <= in_in_update_0_write_write_1_stage_155;
      in_in_update_0_write_write_1_stage_157 <= in_in_update_0_write_write_1_stage_156;
      in_in_update_0_write_write_1_stage_158 <= in_in_update_0_write_write_1_stage_157;
      in_in_update_0_write_write_1_stage_159 <= in_in_update_0_write_write_1_stage_158;
      in_in_update_0_write_write_1_stage_160 <= in_in_update_0_write_write_1_stage_159;
      in_in_update_0_write_write_1_stage_161 <= in_in_update_0_write_write_1_stage_160;
      in_in_update_0_write_write_1_stage_162 <= in_in_update_0_write_write_1_stage_161;
      in_in_update_0_write_write_1_stage_163 <= in_in_update_0_write_write_1_stage_162;
      in_in_update_0_write_write_1_stage_164 <= in_in_update_0_write_write_1_stage_163;
      in_in_update_0_write_write_1_stage_165 <= in_in_update_0_write_write_1_stage_164;
      in_in_update_0_write_write_1_stage_166 <= in_in_update_0_write_write_1_stage_165;
      in_in_update_0_write_write_1_stage_167 <= in_in_update_0_write_write_1_stage_166;
      in_in_update_0_write_write_1_stage_168 <= in_in_update_0_write_write_1_stage_167;
      in_in_update_0_write_write_1_stage_169 <= in_in_update_0_write_write_1_stage_168;
      in_in_update_0_write_write_1_stage_170 <= in_in_update_0_write_write_1_stage_169;
      in_in_update_0_write_write_1_stage_171 <= in_in_update_0_write_write_1_stage_170;
      in_in_update_0_write_write_1_stage_172 <= in_in_update_0_write_write_1_stage_171;
      in_in_update_0_write_write_1_stage_173 <= in_in_update_0_write_write_1_stage_172;
      in_in_update_0_write_write_1_stage_174 <= in_in_update_0_write_write_1_stage_173;
      in_in_update_0_write_write_1_stage_175 <= in_in_update_0_write_write_1_stage_174;
      in_in_update_0_write_write_1_stage_176 <= in_in_update_0_write_write_1_stage_175;
      in_in_update_0_write_write_1_stage_177 <= in_in_update_0_write_write_1_stage_176;
      in_in_update_0_write_write_1_stage_178 <= in_in_update_0_write_write_1_stage_177;
      in_in_update_0_write_write_1_stage_179 <= in_in_update_0_write_write_1_stage_178;
      in_in_update_0_write_write_1_stage_180 <= in_in_update_0_write_write_1_stage_179;
      in_in_update_0_write_write_1_stage_181 <= in_in_update_0_write_write_1_stage_180;
      in_bright_update_0_read_read_2_stage_5 <= in_bright_update_0_read_read_2;
      in_bright_update_0_read_read_2_stage_6 <= in_bright_update_0_read_read_2_stage_5;
      in_bright_update_0_read_read_2_stage_7 <= in_bright_update_0_read_read_2_stage_6;
      in_bright_update_0_read_read_2_stage_8 <= in_bright_update_0_read_read_2_stage_7;
      in_bright_update_0_read_read_2_stage_9 <= in_bright_update_0_read_read_2_stage_8;
      in_bright_update_0_read_read_2_stage_10 <= in_bright_update_0_read_read_2_stage_9;
      in_bright_update_0_read_read_2_stage_11 <= in_bright_update_0_read_read_2_stage_10;
      in_bright_update_0_read_read_2_stage_12 <= in_bright_update_0_read_read_2_stage_11;
      in_bright_update_0_read_read_2_stage_13 <= in_bright_update_0_read_read_2_stage_12;
      in_bright_update_0_read_read_2_stage_14 <= in_bright_update_0_read_read_2_stage_13;
      in_bright_update_0_read_read_2_stage_15 <= in_bright_update_0_read_read_2_stage_14;
      in_bright_update_0_read_read_2_stage_16 <= in_bright_update_0_read_read_2_stage_15;
      in_bright_update_0_read_read_2_stage_17 <= in_bright_update_0_read_read_2_stage_16;
      in_bright_update_0_read_read_2_stage_18 <= in_bright_update_0_read_read_2_stage_17;
      in_bright_update_0_read_read_2_stage_19 <= in_bright_update_0_read_read_2_stage_18;
      in_bright_update_0_read_read_2_stage_20 <= in_bright_update_0_read_read_2_stage_19;
      in_bright_update_0_read_read_2_stage_21 <= in_bright_update_0_read_read_2_stage_20;
      in_bright_update_0_read_read_2_stage_22 <= in_bright_update_0_read_read_2_stage_21;
      in_bright_update_0_read_read_2_stage_23 <= in_bright_update_0_read_read_2_stage_22;
      in_bright_update_0_read_read_2_stage_24 <= in_bright_update_0_read_read_2_stage_23;
      in_bright_update_0_read_read_2_stage_25 <= in_bright_update_0_read_read_2_stage_24;
      in_bright_update_0_read_read_2_stage_26 <= in_bright_update_0_read_read_2_stage_25;
      in_bright_update_0_read_read_2_stage_27 <= in_bright_update_0_read_read_2_stage_26;
      in_bright_update_0_read_read_2_stage_28 <= in_bright_update_0_read_read_2_stage_27;
      in_bright_update_0_read_read_2_stage_29 <= in_bright_update_0_read_read_2_stage_28;
      in_bright_update_0_read_read_2_stage_30 <= in_bright_update_0_read_read_2_stage_29;
      in_bright_update_0_read_read_2_stage_31 <= in_bright_update_0_read_read_2_stage_30;
      in_bright_update_0_read_read_2_stage_32 <= in_bright_update_0_read_read_2_stage_31;
      in_bright_update_0_read_read_2_stage_33 <= in_bright_update_0_read_read_2_stage_32;
      in_bright_update_0_read_read_2_stage_34 <= in_bright_update_0_read_read_2_stage_33;
      in_bright_update_0_read_read_2_stage_35 <= in_bright_update_0_read_read_2_stage_34;
      in_bright_update_0_read_read_2_stage_36 <= in_bright_update_0_read_read_2_stage_35;
      in_bright_update_0_read_read_2_stage_37 <= in_bright_update_0_read_read_2_stage_36;
      in_bright_update_0_read_read_2_stage_38 <= in_bright_update_0_read_read_2_stage_37;
      in_bright_update_0_read_read_2_stage_39 <= in_bright_update_0_read_read_2_stage_38;
      in_bright_update_0_read_read_2_stage_40 <= in_bright_update_0_read_read_2_stage_39;
      in_bright_update_0_read_read_2_stage_41 <= in_bright_update_0_read_read_2_stage_40;
      in_bright_update_0_read_read_2_stage_42 <= in_bright_update_0_read_read_2_stage_41;
      in_bright_update_0_read_read_2_stage_43 <= in_bright_update_0_read_read_2_stage_42;
      in_bright_update_0_read_read_2_stage_44 <= in_bright_update_0_read_read_2_stage_43;
      in_bright_update_0_read_read_2_stage_45 <= in_bright_update_0_read_read_2_stage_44;
      in_bright_update_0_read_read_2_stage_46 <= in_bright_update_0_read_read_2_stage_45;
      in_bright_update_0_read_read_2_stage_47 <= in_bright_update_0_read_read_2_stage_46;
      in_bright_update_0_read_read_2_stage_48 <= in_bright_update_0_read_read_2_stage_47;
      in_bright_update_0_read_read_2_stage_49 <= in_bright_update_0_read_read_2_stage_48;
      in_bright_update_0_read_read_2_stage_50 <= in_bright_update_0_read_read_2_stage_49;
      in_bright_update_0_read_read_2_stage_51 <= in_bright_update_0_read_read_2_stage_50;
      in_bright_update_0_read_read_2_stage_52 <= in_bright_update_0_read_read_2_stage_51;
      in_bright_update_0_read_read_2_stage_53 <= in_bright_update_0_read_read_2_stage_52;
      in_bright_update_0_read_read_2_stage_54 <= in_bright_update_0_read_read_2_stage_53;
      in_bright_update_0_read_read_2_stage_55 <= in_bright_update_0_read_read_2_stage_54;
      in_bright_update_0_read_read_2_stage_56 <= in_bright_update_0_read_read_2_stage_55;
      in_bright_update_0_read_read_2_stage_57 <= in_bright_update_0_read_read_2_stage_56;
      in_bright_update_0_read_read_2_stage_58 <= in_bright_update_0_read_read_2_stage_57;
      in_bright_update_0_read_read_2_stage_59 <= in_bright_update_0_read_read_2_stage_58;
      in_bright_update_0_read_read_2_stage_60 <= in_bright_update_0_read_read_2_stage_59;
      in_bright_update_0_read_read_2_stage_61 <= in_bright_update_0_read_read_2_stage_60;
      in_bright_update_0_read_read_2_stage_62 <= in_bright_update_0_read_read_2_stage_61;
      in_bright_update_0_read_read_2_stage_63 <= in_bright_update_0_read_read_2_stage_62;
      in_bright_update_0_read_read_2_stage_64 <= in_bright_update_0_read_read_2_stage_63;
      in_bright_update_0_read_read_2_stage_65 <= in_bright_update_0_read_read_2_stage_64;
      in_bright_update_0_read_read_2_stage_66 <= in_bright_update_0_read_read_2_stage_65;
      in_bright_update_0_read_read_2_stage_67 <= in_bright_update_0_read_read_2_stage_66;
      in_bright_update_0_read_read_2_stage_68 <= in_bright_update_0_read_read_2_stage_67;
      in_bright_update_0_read_read_2_stage_69 <= in_bright_update_0_read_read_2_stage_68;
      in_bright_update_0_read_read_2_stage_70 <= in_bright_update_0_read_read_2_stage_69;
      in_bright_update_0_read_read_2_stage_71 <= in_bright_update_0_read_read_2_stage_70;
      in_bright_update_0_read_read_2_stage_72 <= in_bright_update_0_read_read_2_stage_71;
      in_bright_update_0_read_read_2_stage_73 <= in_bright_update_0_read_read_2_stage_72;
      in_bright_update_0_read_read_2_stage_74 <= in_bright_update_0_read_read_2_stage_73;
      in_bright_update_0_read_read_2_stage_75 <= in_bright_update_0_read_read_2_stage_74;
      in_bright_update_0_read_read_2_stage_76 <= in_bright_update_0_read_read_2_stage_75;
      in_bright_update_0_read_read_2_stage_77 <= in_bright_update_0_read_read_2_stage_76;
      in_bright_update_0_read_read_2_stage_78 <= in_bright_update_0_read_read_2_stage_77;
      in_bright_update_0_read_read_2_stage_79 <= in_bright_update_0_read_read_2_stage_78;
      in_bright_update_0_read_read_2_stage_80 <= in_bright_update_0_read_read_2_stage_79;
      in_bright_update_0_read_read_2_stage_81 <= in_bright_update_0_read_read_2_stage_80;
      in_bright_update_0_read_read_2_stage_82 <= in_bright_update_0_read_read_2_stage_81;
      in_bright_update_0_read_read_2_stage_83 <= in_bright_update_0_read_read_2_stage_82;
      in_bright_update_0_read_read_2_stage_84 <= in_bright_update_0_read_read_2_stage_83;
      in_bright_update_0_read_read_2_stage_85 <= in_bright_update_0_read_read_2_stage_84;
      in_bright_update_0_read_read_2_stage_86 <= in_bright_update_0_read_read_2_stage_85;
      in_bright_update_0_read_read_2_stage_87 <= in_bright_update_0_read_read_2_stage_86;
      in_bright_update_0_read_read_2_stage_88 <= in_bright_update_0_read_read_2_stage_87;
      in_bright_update_0_read_read_2_stage_89 <= in_bright_update_0_read_read_2_stage_88;
      in_bright_update_0_read_read_2_stage_90 <= in_bright_update_0_read_read_2_stage_89;
      in_bright_update_0_read_read_2_stage_91 <= in_bright_update_0_read_read_2_stage_90;
      in_bright_update_0_read_read_2_stage_92 <= in_bright_update_0_read_read_2_stage_91;
      in_bright_update_0_read_read_2_stage_93 <= in_bright_update_0_read_read_2_stage_92;
      in_bright_update_0_read_read_2_stage_94 <= in_bright_update_0_read_read_2_stage_93;
      in_bright_update_0_read_read_2_stage_95 <= in_bright_update_0_read_read_2_stage_94;
      in_bright_update_0_read_read_2_stage_96 <= in_bright_update_0_read_read_2_stage_95;
      in_bright_update_0_read_read_2_stage_97 <= in_bright_update_0_read_read_2_stage_96;
      in_bright_update_0_read_read_2_stage_98 <= in_bright_update_0_read_read_2_stage_97;
      in_bright_update_0_read_read_2_stage_99 <= in_bright_update_0_read_read_2_stage_98;
      in_bright_update_0_read_read_2_stage_100 <= in_bright_update_0_read_read_2_stage_99;
      in_bright_update_0_read_read_2_stage_101 <= in_bright_update_0_read_read_2_stage_100;
      in_bright_update_0_read_read_2_stage_102 <= in_bright_update_0_read_read_2_stage_101;
      in_bright_update_0_read_read_2_stage_103 <= in_bright_update_0_read_read_2_stage_102;
      in_bright_update_0_read_read_2_stage_104 <= in_bright_update_0_read_read_2_stage_103;
      in_bright_update_0_read_read_2_stage_105 <= in_bright_update_0_read_read_2_stage_104;
      in_bright_update_0_read_read_2_stage_106 <= in_bright_update_0_read_read_2_stage_105;
      in_bright_update_0_read_read_2_stage_107 <= in_bright_update_0_read_read_2_stage_106;
      in_bright_update_0_read_read_2_stage_108 <= in_bright_update_0_read_read_2_stage_107;
      in_bright_update_0_read_read_2_stage_109 <= in_bright_update_0_read_read_2_stage_108;
      in_bright_update_0_read_read_2_stage_110 <= in_bright_update_0_read_read_2_stage_109;
      in_bright_update_0_read_read_2_stage_111 <= in_bright_update_0_read_read_2_stage_110;
      in_bright_update_0_read_read_2_stage_112 <= in_bright_update_0_read_read_2_stage_111;
      in_bright_update_0_read_read_2_stage_113 <= in_bright_update_0_read_read_2_stage_112;
      in_bright_update_0_read_read_2_stage_114 <= in_bright_update_0_read_read_2_stage_113;
      in_bright_update_0_read_read_2_stage_115 <= in_bright_update_0_read_read_2_stage_114;
      in_bright_update_0_read_read_2_stage_116 <= in_bright_update_0_read_read_2_stage_115;
      in_bright_update_0_read_read_2_stage_117 <= in_bright_update_0_read_read_2_stage_116;
      in_bright_update_0_read_read_2_stage_118 <= in_bright_update_0_read_read_2_stage_117;
      in_bright_update_0_read_read_2_stage_119 <= in_bright_update_0_read_read_2_stage_118;
      in_bright_update_0_read_read_2_stage_120 <= in_bright_update_0_read_read_2_stage_119;
      in_bright_update_0_read_read_2_stage_121 <= in_bright_update_0_read_read_2_stage_120;
      in_bright_update_0_read_read_2_stage_122 <= in_bright_update_0_read_read_2_stage_121;
      in_bright_update_0_read_read_2_stage_123 <= in_bright_update_0_read_read_2_stage_122;
      in_bright_update_0_read_read_2_stage_124 <= in_bright_update_0_read_read_2_stage_123;
      in_bright_update_0_read_read_2_stage_125 <= in_bright_update_0_read_read_2_stage_124;
      in_bright_update_0_read_read_2_stage_126 <= in_bright_update_0_read_read_2_stage_125;
      in_bright_update_0_read_read_2_stage_127 <= in_bright_update_0_read_read_2_stage_126;
      in_bright_update_0_read_read_2_stage_128 <= in_bright_update_0_read_read_2_stage_127;
      in_bright_update_0_read_read_2_stage_129 <= in_bright_update_0_read_read_2_stage_128;
      in_bright_update_0_read_read_2_stage_130 <= in_bright_update_0_read_read_2_stage_129;
      in_bright_update_0_read_read_2_stage_131 <= in_bright_update_0_read_read_2_stage_130;
      in_bright_update_0_read_read_2_stage_132 <= in_bright_update_0_read_read_2_stage_131;
      in_bright_update_0_read_read_2_stage_133 <= in_bright_update_0_read_read_2_stage_132;
      in_bright_update_0_read_read_2_stage_134 <= in_bright_update_0_read_read_2_stage_133;
      in_bright_update_0_read_read_2_stage_135 <= in_bright_update_0_read_read_2_stage_134;
      in_bright_update_0_read_read_2_stage_136 <= in_bright_update_0_read_read_2_stage_135;
      in_bright_update_0_read_read_2_stage_137 <= in_bright_update_0_read_read_2_stage_136;
      in_bright_update_0_read_read_2_stage_138 <= in_bright_update_0_read_read_2_stage_137;
      in_bright_update_0_read_read_2_stage_139 <= in_bright_update_0_read_read_2_stage_138;
      in_bright_update_0_read_read_2_stage_140 <= in_bright_update_0_read_read_2_stage_139;
      in_bright_update_0_read_read_2_stage_141 <= in_bright_update_0_read_read_2_stage_140;
      in_bright_update_0_read_read_2_stage_142 <= in_bright_update_0_read_read_2_stage_141;
      in_bright_update_0_read_read_2_stage_143 <= in_bright_update_0_read_read_2_stage_142;
      in_bright_update_0_read_read_2_stage_144 <= in_bright_update_0_read_read_2_stage_143;
      in_bright_update_0_read_read_2_stage_145 <= in_bright_update_0_read_read_2_stage_144;
      in_bright_update_0_read_read_2_stage_146 <= in_bright_update_0_read_read_2_stage_145;
      in_bright_update_0_read_read_2_stage_147 <= in_bright_update_0_read_read_2_stage_146;
      in_bright_update_0_read_read_2_stage_148 <= in_bright_update_0_read_read_2_stage_147;
      in_bright_update_0_read_read_2_stage_149 <= in_bright_update_0_read_read_2_stage_148;
      in_bright_update_0_read_read_2_stage_150 <= in_bright_update_0_read_read_2_stage_149;
      in_bright_update_0_read_read_2_stage_151 <= in_bright_update_0_read_read_2_stage_150;
      in_bright_update_0_read_read_2_stage_152 <= in_bright_update_0_read_read_2_stage_151;
      in_bright_update_0_read_read_2_stage_153 <= in_bright_update_0_read_read_2_stage_152;
      in_bright_update_0_read_read_2_stage_154 <= in_bright_update_0_read_read_2_stage_153;
      in_bright_update_0_read_read_2_stage_155 <= in_bright_update_0_read_read_2_stage_154;
      in_bright_update_0_read_read_2_stage_156 <= in_bright_update_0_read_read_2_stage_155;
      in_bright_update_0_read_read_2_stage_157 <= in_bright_update_0_read_read_2_stage_156;
      in_bright_update_0_read_read_2_stage_158 <= in_bright_update_0_read_read_2_stage_157;
      in_bright_update_0_read_read_2_stage_159 <= in_bright_update_0_read_read_2_stage_158;
      in_bright_update_0_read_read_2_stage_160 <= in_bright_update_0_read_read_2_stage_159;
      in_bright_update_0_read_read_2_stage_161 <= in_bright_update_0_read_read_2_stage_160;
      in_bright_update_0_read_read_2_stage_162 <= in_bright_update_0_read_read_2_stage_161;
      in_bright_update_0_read_read_2_stage_163 <= in_bright_update_0_read_read_2_stage_162;
      in_bright_update_0_read_read_2_stage_164 <= in_bright_update_0_read_read_2_stage_163;
      in_bright_update_0_read_read_2_stage_165 <= in_bright_update_0_read_read_2_stage_164;
      in_bright_update_0_read_read_2_stage_166 <= in_bright_update_0_read_read_2_stage_165;
      in_bright_update_0_read_read_2_stage_167 <= in_bright_update_0_read_read_2_stage_166;
      in_bright_update_0_read_read_2_stage_168 <= in_bright_update_0_read_read_2_stage_167;
      in_bright_update_0_read_read_2_stage_169 <= in_bright_update_0_read_read_2_stage_168;
      in_bright_update_0_read_read_2_stage_170 <= in_bright_update_0_read_read_2_stage_169;
      in_bright_update_0_read_read_2_stage_171 <= in_bright_update_0_read_read_2_stage_170;
      in_bright_update_0_read_read_2_stage_172 <= in_bright_update_0_read_read_2_stage_171;
      in_bright_update_0_read_read_2_stage_173 <= in_bright_update_0_read_read_2_stage_172;
      in_bright_update_0_read_read_2_stage_174 <= in_bright_update_0_read_read_2_stage_173;
      in_bright_update_0_read_read_2_stage_175 <= in_bright_update_0_read_read_2_stage_174;
      in_bright_update_0_read_read_2_stage_176 <= in_bright_update_0_read_read_2_stage_175;
      in_bright_update_0_read_read_2_stage_177 <= in_bright_update_0_read_read_2_stage_176;
      in_bright_update_0_read_read_2_stage_178 <= in_bright_update_0_read_read_2_stage_177;
      in_bright_update_0_read_read_2_stage_179 <= in_bright_update_0_read_read_2_stage_178;
      in_bright_update_0_read_read_2_stage_180 <= in_bright_update_0_read_read_2_stage_179;
      in_bright_update_0_read_read_2_stage_181 <= in_bright_update_0_read_read_2_stage_180;
      bright_update_0_stage_6 <= bright_update_0;
      bright_update_0_stage_7 <= bright_update_0_stage_6;
      bright_update_0_stage_8 <= bright_update_0_stage_7;
      bright_update_0_stage_9 <= bright_update_0_stage_8;
      bright_update_0_stage_10 <= bright_update_0_stage_9;
      bright_update_0_stage_11 <= bright_update_0_stage_10;
      bright_update_0_stage_12 <= bright_update_0_stage_11;
      bright_update_0_stage_13 <= bright_update_0_stage_12;
      bright_update_0_stage_14 <= bright_update_0_stage_13;
      bright_update_0_stage_15 <= bright_update_0_stage_14;
      bright_update_0_stage_16 <= bright_update_0_stage_15;
      bright_update_0_stage_17 <= bright_update_0_stage_16;
      bright_update_0_stage_18 <= bright_update_0_stage_17;
      bright_update_0_stage_19 <= bright_update_0_stage_18;
      bright_update_0_stage_20 <= bright_update_0_stage_19;
      bright_update_0_stage_21 <= bright_update_0_stage_20;
      bright_update_0_stage_22 <= bright_update_0_stage_21;
      bright_update_0_stage_23 <= bright_update_0_stage_22;
      bright_update_0_stage_24 <= bright_update_0_stage_23;
      bright_update_0_stage_25 <= bright_update_0_stage_24;
      bright_update_0_stage_26 <= bright_update_0_stage_25;
      bright_update_0_stage_27 <= bright_update_0_stage_26;
      bright_update_0_stage_28 <= bright_update_0_stage_27;
      bright_update_0_stage_29 <= bright_update_0_stage_28;
      bright_update_0_stage_30 <= bright_update_0_stage_29;
      bright_update_0_stage_31 <= bright_update_0_stage_30;
      bright_update_0_stage_32 <= bright_update_0_stage_31;
      bright_update_0_stage_33 <= bright_update_0_stage_32;
      bright_update_0_stage_34 <= bright_update_0_stage_33;
      bright_update_0_stage_35 <= bright_update_0_stage_34;
      bright_update_0_stage_36 <= bright_update_0_stage_35;
      bright_update_0_stage_37 <= bright_update_0_stage_36;
      bright_update_0_stage_38 <= bright_update_0_stage_37;
      bright_update_0_stage_39 <= bright_update_0_stage_38;
      bright_update_0_stage_40 <= bright_update_0_stage_39;
      bright_update_0_stage_41 <= bright_update_0_stage_40;
      bright_update_0_stage_42 <= bright_update_0_stage_41;
      bright_update_0_stage_43 <= bright_update_0_stage_42;
      bright_update_0_stage_44 <= bright_update_0_stage_43;
      bright_update_0_stage_45 <= bright_update_0_stage_44;
      bright_update_0_stage_46 <= bright_update_0_stage_45;
      bright_update_0_stage_47 <= bright_update_0_stage_46;
      bright_update_0_stage_48 <= bright_update_0_stage_47;
      bright_update_0_stage_49 <= bright_update_0_stage_48;
      bright_update_0_stage_50 <= bright_update_0_stage_49;
      bright_update_0_stage_51 <= bright_update_0_stage_50;
      bright_update_0_stage_52 <= bright_update_0_stage_51;
      bright_update_0_stage_53 <= bright_update_0_stage_52;
      bright_update_0_stage_54 <= bright_update_0_stage_53;
      bright_update_0_stage_55 <= bright_update_0_stage_54;
      bright_update_0_stage_56 <= bright_update_0_stage_55;
      bright_update_0_stage_57 <= bright_update_0_stage_56;
      bright_update_0_stage_58 <= bright_update_0_stage_57;
      bright_update_0_stage_59 <= bright_update_0_stage_58;
      bright_update_0_stage_60 <= bright_update_0_stage_59;
      bright_update_0_stage_61 <= bright_update_0_stage_60;
      bright_update_0_stage_62 <= bright_update_0_stage_61;
      bright_update_0_stage_63 <= bright_update_0_stage_62;
      bright_update_0_stage_64 <= bright_update_0_stage_63;
      bright_update_0_stage_65 <= bright_update_0_stage_64;
      bright_update_0_stage_66 <= bright_update_0_stage_65;
      bright_update_0_stage_67 <= bright_update_0_stage_66;
      bright_update_0_stage_68 <= bright_update_0_stage_67;
      bright_update_0_stage_69 <= bright_update_0_stage_68;
      bright_update_0_stage_70 <= bright_update_0_stage_69;
      bright_update_0_stage_71 <= bright_update_0_stage_70;
      bright_update_0_stage_72 <= bright_update_0_stage_71;
      bright_update_0_stage_73 <= bright_update_0_stage_72;
      bright_update_0_stage_74 <= bright_update_0_stage_73;
      bright_update_0_stage_75 <= bright_update_0_stage_74;
      bright_update_0_stage_76 <= bright_update_0_stage_75;
      bright_update_0_stage_77 <= bright_update_0_stage_76;
      bright_update_0_stage_78 <= bright_update_0_stage_77;
      bright_update_0_stage_79 <= bright_update_0_stage_78;
      bright_update_0_stage_80 <= bright_update_0_stage_79;
      bright_update_0_stage_81 <= bright_update_0_stage_80;
      bright_update_0_stage_82 <= bright_update_0_stage_81;
      bright_update_0_stage_83 <= bright_update_0_stage_82;
      bright_update_0_stage_84 <= bright_update_0_stage_83;
      bright_update_0_stage_85 <= bright_update_0_stage_84;
      bright_update_0_stage_86 <= bright_update_0_stage_85;
      bright_update_0_stage_87 <= bright_update_0_stage_86;
      bright_update_0_stage_88 <= bright_update_0_stage_87;
      bright_update_0_stage_89 <= bright_update_0_stage_88;
      bright_update_0_stage_90 <= bright_update_0_stage_89;
      bright_update_0_stage_91 <= bright_update_0_stage_90;
      bright_update_0_stage_92 <= bright_update_0_stage_91;
      bright_update_0_stage_93 <= bright_update_0_stage_92;
      bright_update_0_stage_94 <= bright_update_0_stage_93;
      bright_update_0_stage_95 <= bright_update_0_stage_94;
      bright_update_0_stage_96 <= bright_update_0_stage_95;
      bright_update_0_stage_97 <= bright_update_0_stage_96;
      bright_update_0_stage_98 <= bright_update_0_stage_97;
      bright_update_0_stage_99 <= bright_update_0_stage_98;
      bright_update_0_stage_100 <= bright_update_0_stage_99;
      bright_update_0_stage_101 <= bright_update_0_stage_100;
      bright_update_0_stage_102 <= bright_update_0_stage_101;
      bright_update_0_stage_103 <= bright_update_0_stage_102;
      bright_update_0_stage_104 <= bright_update_0_stage_103;
      bright_update_0_stage_105 <= bright_update_0_stage_104;
      bright_update_0_stage_106 <= bright_update_0_stage_105;
      bright_update_0_stage_107 <= bright_update_0_stage_106;
      bright_update_0_stage_108 <= bright_update_0_stage_107;
      bright_update_0_stage_109 <= bright_update_0_stage_108;
      bright_update_0_stage_110 <= bright_update_0_stage_109;
      bright_update_0_stage_111 <= bright_update_0_stage_110;
      bright_update_0_stage_112 <= bright_update_0_stage_111;
      bright_update_0_stage_113 <= bright_update_0_stage_112;
      bright_update_0_stage_114 <= bright_update_0_stage_113;
      bright_update_0_stage_115 <= bright_update_0_stage_114;
      bright_update_0_stage_116 <= bright_update_0_stage_115;
      bright_update_0_stage_117 <= bright_update_0_stage_116;
      bright_update_0_stage_118 <= bright_update_0_stage_117;
      bright_update_0_stage_119 <= bright_update_0_stage_118;
      bright_update_0_stage_120 <= bright_update_0_stage_119;
      bright_update_0_stage_121 <= bright_update_0_stage_120;
      bright_update_0_stage_122 <= bright_update_0_stage_121;
      bright_update_0_stage_123 <= bright_update_0_stage_122;
      bright_update_0_stage_124 <= bright_update_0_stage_123;
      bright_update_0_stage_125 <= bright_update_0_stage_124;
      bright_update_0_stage_126 <= bright_update_0_stage_125;
      bright_update_0_stage_127 <= bright_update_0_stage_126;
      bright_update_0_stage_128 <= bright_update_0_stage_127;
      bright_update_0_stage_129 <= bright_update_0_stage_128;
      bright_update_0_stage_130 <= bright_update_0_stage_129;
      bright_update_0_stage_131 <= bright_update_0_stage_130;
      bright_update_0_stage_132 <= bright_update_0_stage_131;
      bright_update_0_stage_133 <= bright_update_0_stage_132;
      bright_update_0_stage_134 <= bright_update_0_stage_133;
      bright_update_0_stage_135 <= bright_update_0_stage_134;
      bright_update_0_stage_136 <= bright_update_0_stage_135;
      bright_update_0_stage_137 <= bright_update_0_stage_136;
      bright_update_0_stage_138 <= bright_update_0_stage_137;
      bright_update_0_stage_139 <= bright_update_0_stage_138;
      bright_update_0_stage_140 <= bright_update_0_stage_139;
      bright_update_0_stage_141 <= bright_update_0_stage_140;
      bright_update_0_stage_142 <= bright_update_0_stage_141;
      bright_update_0_stage_143 <= bright_update_0_stage_142;
      bright_update_0_stage_144 <= bright_update_0_stage_143;
      bright_update_0_stage_145 <= bright_update_0_stage_144;
      bright_update_0_stage_146 <= bright_update_0_stage_145;
      bright_update_0_stage_147 <= bright_update_0_stage_146;
      bright_update_0_stage_148 <= bright_update_0_stage_147;
      bright_update_0_stage_149 <= bright_update_0_stage_148;
      bright_update_0_stage_150 <= bright_update_0_stage_149;
      bright_update_0_stage_151 <= bright_update_0_stage_150;
      bright_update_0_stage_152 <= bright_update_0_stage_151;
      bright_update_0_stage_153 <= bright_update_0_stage_152;
      bright_update_0_stage_154 <= bright_update_0_stage_153;
      bright_update_0_stage_155 <= bright_update_0_stage_154;
      bright_update_0_stage_156 <= bright_update_0_stage_155;
      bright_update_0_stage_157 <= bright_update_0_stage_156;
      bright_update_0_stage_158 <= bright_update_0_stage_157;
      bright_update_0_stage_159 <= bright_update_0_stage_158;
      bright_update_0_stage_160 <= bright_update_0_stage_159;
      bright_update_0_stage_161 <= bright_update_0_stage_160;
      bright_update_0_stage_162 <= bright_update_0_stage_161;
      bright_update_0_stage_163 <= bright_update_0_stage_162;
      bright_update_0_stage_164 <= bright_update_0_stage_163;
      bright_update_0_stage_165 <= bright_update_0_stage_164;
      bright_update_0_stage_166 <= bright_update_0_stage_165;
      bright_update_0_stage_167 <= bright_update_0_stage_166;
      bright_update_0_stage_168 <= bright_update_0_stage_167;
      bright_update_0_stage_169 <= bright_update_0_stage_168;
      bright_update_0_stage_170 <= bright_update_0_stage_169;
      bright_update_0_stage_171 <= bright_update_0_stage_170;
      bright_update_0_stage_172 <= bright_update_0_stage_171;
      bright_update_0_stage_173 <= bright_update_0_stage_172;
      bright_update_0_stage_174 <= bright_update_0_stage_173;
      bright_update_0_stage_175 <= bright_update_0_stage_174;
      bright_update_0_stage_176 <= bright_update_0_stage_175;
      bright_update_0_stage_177 <= bright_update_0_stage_176;
      bright_update_0_stage_178 <= bright_update_0_stage_177;
      bright_update_0_stage_179 <= bright_update_0_stage_178;
      bright_update_0_stage_180 <= bright_update_0_stage_179;
      bright_update_0_stage_181 <= bright_update_0_stage_180;
      bright_bright_update_0_write_write_3_stage_7 <= bright_bright_update_0_write_write_3;
      bright_bright_update_0_write_write_3_stage_8 <= bright_bright_update_0_write_write_3_stage_7;
      bright_bright_update_0_write_write_3_stage_9 <= bright_bright_update_0_write_write_3_stage_8;
      bright_bright_update_0_write_write_3_stage_10 <= bright_bright_update_0_write_write_3_stage_9;
      bright_bright_update_0_write_write_3_stage_11 <= bright_bright_update_0_write_write_3_stage_10;
      bright_bright_update_0_write_write_3_stage_12 <= bright_bright_update_0_write_write_3_stage_11;
      bright_bright_update_0_write_write_3_stage_13 <= bright_bright_update_0_write_write_3_stage_12;
      bright_bright_update_0_write_write_3_stage_14 <= bright_bright_update_0_write_write_3_stage_13;
      bright_bright_update_0_write_write_3_stage_15 <= bright_bright_update_0_write_write_3_stage_14;
      bright_bright_update_0_write_write_3_stage_16 <= bright_bright_update_0_write_write_3_stage_15;
      bright_bright_update_0_write_write_3_stage_17 <= bright_bright_update_0_write_write_3_stage_16;
      bright_bright_update_0_write_write_3_stage_18 <= bright_bright_update_0_write_write_3_stage_17;
      bright_bright_update_0_write_write_3_stage_19 <= bright_bright_update_0_write_write_3_stage_18;
      bright_bright_update_0_write_write_3_stage_20 <= bright_bright_update_0_write_write_3_stage_19;
      bright_bright_update_0_write_write_3_stage_21 <= bright_bright_update_0_write_write_3_stage_20;
      bright_bright_update_0_write_write_3_stage_22 <= bright_bright_update_0_write_write_3_stage_21;
      bright_bright_update_0_write_write_3_stage_23 <= bright_bright_update_0_write_write_3_stage_22;
      bright_bright_update_0_write_write_3_stage_24 <= bright_bright_update_0_write_write_3_stage_23;
      bright_bright_update_0_write_write_3_stage_25 <= bright_bright_update_0_write_write_3_stage_24;
      bright_bright_update_0_write_write_3_stage_26 <= bright_bright_update_0_write_write_3_stage_25;
      bright_bright_update_0_write_write_3_stage_27 <= bright_bright_update_0_write_write_3_stage_26;
      bright_bright_update_0_write_write_3_stage_28 <= bright_bright_update_0_write_write_3_stage_27;
      bright_bright_update_0_write_write_3_stage_29 <= bright_bright_update_0_write_write_3_stage_28;
      bright_bright_update_0_write_write_3_stage_30 <= bright_bright_update_0_write_write_3_stage_29;
      bright_bright_update_0_write_write_3_stage_31 <= bright_bright_update_0_write_write_3_stage_30;
      bright_bright_update_0_write_write_3_stage_32 <= bright_bright_update_0_write_write_3_stage_31;
      bright_bright_update_0_write_write_3_stage_33 <= bright_bright_update_0_write_write_3_stage_32;
      bright_bright_update_0_write_write_3_stage_34 <= bright_bright_update_0_write_write_3_stage_33;
      bright_bright_update_0_write_write_3_stage_35 <= bright_bright_update_0_write_write_3_stage_34;
      bright_bright_update_0_write_write_3_stage_36 <= bright_bright_update_0_write_write_3_stage_35;
      bright_bright_update_0_write_write_3_stage_37 <= bright_bright_update_0_write_write_3_stage_36;
      bright_bright_update_0_write_write_3_stage_38 <= bright_bright_update_0_write_write_3_stage_37;
      bright_bright_update_0_write_write_3_stage_39 <= bright_bright_update_0_write_write_3_stage_38;
      bright_bright_update_0_write_write_3_stage_40 <= bright_bright_update_0_write_write_3_stage_39;
      bright_bright_update_0_write_write_3_stage_41 <= bright_bright_update_0_write_write_3_stage_40;
      bright_bright_update_0_write_write_3_stage_42 <= bright_bright_update_0_write_write_3_stage_41;
      bright_bright_update_0_write_write_3_stage_43 <= bright_bright_update_0_write_write_3_stage_42;
      bright_bright_update_0_write_write_3_stage_44 <= bright_bright_update_0_write_write_3_stage_43;
      bright_bright_update_0_write_write_3_stage_45 <= bright_bright_update_0_write_write_3_stage_44;
      bright_bright_update_0_write_write_3_stage_46 <= bright_bright_update_0_write_write_3_stage_45;
      bright_bright_update_0_write_write_3_stage_47 <= bright_bright_update_0_write_write_3_stage_46;
      bright_bright_update_0_write_write_3_stage_48 <= bright_bright_update_0_write_write_3_stage_47;
      bright_bright_update_0_write_write_3_stage_49 <= bright_bright_update_0_write_write_3_stage_48;
      bright_bright_update_0_write_write_3_stage_50 <= bright_bright_update_0_write_write_3_stage_49;
      bright_bright_update_0_write_write_3_stage_51 <= bright_bright_update_0_write_write_3_stage_50;
      bright_bright_update_0_write_write_3_stage_52 <= bright_bright_update_0_write_write_3_stage_51;
      bright_bright_update_0_write_write_3_stage_53 <= bright_bright_update_0_write_write_3_stage_52;
      bright_bright_update_0_write_write_3_stage_54 <= bright_bright_update_0_write_write_3_stage_53;
      bright_bright_update_0_write_write_3_stage_55 <= bright_bright_update_0_write_write_3_stage_54;
      bright_bright_update_0_write_write_3_stage_56 <= bright_bright_update_0_write_write_3_stage_55;
      bright_bright_update_0_write_write_3_stage_57 <= bright_bright_update_0_write_write_3_stage_56;
      bright_bright_update_0_write_write_3_stage_58 <= bright_bright_update_0_write_write_3_stage_57;
      bright_bright_update_0_write_write_3_stage_59 <= bright_bright_update_0_write_write_3_stage_58;
      bright_bright_update_0_write_write_3_stage_60 <= bright_bright_update_0_write_write_3_stage_59;
      bright_bright_update_0_write_write_3_stage_61 <= bright_bright_update_0_write_write_3_stage_60;
      bright_bright_update_0_write_write_3_stage_62 <= bright_bright_update_0_write_write_3_stage_61;
      bright_bright_update_0_write_write_3_stage_63 <= bright_bright_update_0_write_write_3_stage_62;
      bright_bright_update_0_write_write_3_stage_64 <= bright_bright_update_0_write_write_3_stage_63;
      bright_bright_update_0_write_write_3_stage_65 <= bright_bright_update_0_write_write_3_stage_64;
      bright_bright_update_0_write_write_3_stage_66 <= bright_bright_update_0_write_write_3_stage_65;
      bright_bright_update_0_write_write_3_stage_67 <= bright_bright_update_0_write_write_3_stage_66;
      bright_bright_update_0_write_write_3_stage_68 <= bright_bright_update_0_write_write_3_stage_67;
      bright_bright_update_0_write_write_3_stage_69 <= bright_bright_update_0_write_write_3_stage_68;
      bright_bright_update_0_write_write_3_stage_70 <= bright_bright_update_0_write_write_3_stage_69;
      bright_bright_update_0_write_write_3_stage_71 <= bright_bright_update_0_write_write_3_stage_70;
      bright_bright_update_0_write_write_3_stage_72 <= bright_bright_update_0_write_write_3_stage_71;
      bright_bright_update_0_write_write_3_stage_73 <= bright_bright_update_0_write_write_3_stage_72;
      bright_bright_update_0_write_write_3_stage_74 <= bright_bright_update_0_write_write_3_stage_73;
      bright_bright_update_0_write_write_3_stage_75 <= bright_bright_update_0_write_write_3_stage_74;
      bright_bright_update_0_write_write_3_stage_76 <= bright_bright_update_0_write_write_3_stage_75;
      bright_bright_update_0_write_write_3_stage_77 <= bright_bright_update_0_write_write_3_stage_76;
      bright_bright_update_0_write_write_3_stage_78 <= bright_bright_update_0_write_write_3_stage_77;
      bright_bright_update_0_write_write_3_stage_79 <= bright_bright_update_0_write_write_3_stage_78;
      bright_bright_update_0_write_write_3_stage_80 <= bright_bright_update_0_write_write_3_stage_79;
      bright_bright_update_0_write_write_3_stage_81 <= bright_bright_update_0_write_write_3_stage_80;
      bright_bright_update_0_write_write_3_stage_82 <= bright_bright_update_0_write_write_3_stage_81;
      bright_bright_update_0_write_write_3_stage_83 <= bright_bright_update_0_write_write_3_stage_82;
      bright_bright_update_0_write_write_3_stage_84 <= bright_bright_update_0_write_write_3_stage_83;
      bright_bright_update_0_write_write_3_stage_85 <= bright_bright_update_0_write_write_3_stage_84;
      bright_bright_update_0_write_write_3_stage_86 <= bright_bright_update_0_write_write_3_stage_85;
      bright_bright_update_0_write_write_3_stage_87 <= bright_bright_update_0_write_write_3_stage_86;
      bright_bright_update_0_write_write_3_stage_88 <= bright_bright_update_0_write_write_3_stage_87;
      bright_bright_update_0_write_write_3_stage_89 <= bright_bright_update_0_write_write_3_stage_88;
      bright_bright_update_0_write_write_3_stage_90 <= bright_bright_update_0_write_write_3_stage_89;
      bright_bright_update_0_write_write_3_stage_91 <= bright_bright_update_0_write_write_3_stage_90;
      bright_bright_update_0_write_write_3_stage_92 <= bright_bright_update_0_write_write_3_stage_91;
      bright_bright_update_0_write_write_3_stage_93 <= bright_bright_update_0_write_write_3_stage_92;
      bright_bright_update_0_write_write_3_stage_94 <= bright_bright_update_0_write_write_3_stage_93;
      bright_bright_update_0_write_write_3_stage_95 <= bright_bright_update_0_write_write_3_stage_94;
      bright_bright_update_0_write_write_3_stage_96 <= bright_bright_update_0_write_write_3_stage_95;
      bright_bright_update_0_write_write_3_stage_97 <= bright_bright_update_0_write_write_3_stage_96;
      bright_bright_update_0_write_write_3_stage_98 <= bright_bright_update_0_write_write_3_stage_97;
      bright_bright_update_0_write_write_3_stage_99 <= bright_bright_update_0_write_write_3_stage_98;
      bright_bright_update_0_write_write_3_stage_100 <= bright_bright_update_0_write_write_3_stage_99;
      bright_bright_update_0_write_write_3_stage_101 <= bright_bright_update_0_write_write_3_stage_100;
      bright_bright_update_0_write_write_3_stage_102 <= bright_bright_update_0_write_write_3_stage_101;
      bright_bright_update_0_write_write_3_stage_103 <= bright_bright_update_0_write_write_3_stage_102;
      bright_bright_update_0_write_write_3_stage_104 <= bright_bright_update_0_write_write_3_stage_103;
      bright_bright_update_0_write_write_3_stage_105 <= bright_bright_update_0_write_write_3_stage_104;
      bright_bright_update_0_write_write_3_stage_106 <= bright_bright_update_0_write_write_3_stage_105;
      bright_bright_update_0_write_write_3_stage_107 <= bright_bright_update_0_write_write_3_stage_106;
      bright_bright_update_0_write_write_3_stage_108 <= bright_bright_update_0_write_write_3_stage_107;
      bright_bright_update_0_write_write_3_stage_109 <= bright_bright_update_0_write_write_3_stage_108;
      bright_bright_update_0_write_write_3_stage_110 <= bright_bright_update_0_write_write_3_stage_109;
      bright_bright_update_0_write_write_3_stage_111 <= bright_bright_update_0_write_write_3_stage_110;
      bright_bright_update_0_write_write_3_stage_112 <= bright_bright_update_0_write_write_3_stage_111;
      bright_bright_update_0_write_write_3_stage_113 <= bright_bright_update_0_write_write_3_stage_112;
      bright_bright_update_0_write_write_3_stage_114 <= bright_bright_update_0_write_write_3_stage_113;
      bright_bright_update_0_write_write_3_stage_115 <= bright_bright_update_0_write_write_3_stage_114;
      bright_bright_update_0_write_write_3_stage_116 <= bright_bright_update_0_write_write_3_stage_115;
      bright_bright_update_0_write_write_3_stage_117 <= bright_bright_update_0_write_write_3_stage_116;
      bright_bright_update_0_write_write_3_stage_118 <= bright_bright_update_0_write_write_3_stage_117;
      bright_bright_update_0_write_write_3_stage_119 <= bright_bright_update_0_write_write_3_stage_118;
      bright_bright_update_0_write_write_3_stage_120 <= bright_bright_update_0_write_write_3_stage_119;
      bright_bright_update_0_write_write_3_stage_121 <= bright_bright_update_0_write_write_3_stage_120;
      bright_bright_update_0_write_write_3_stage_122 <= bright_bright_update_0_write_write_3_stage_121;
      bright_bright_update_0_write_write_3_stage_123 <= bright_bright_update_0_write_write_3_stage_122;
      bright_bright_update_0_write_write_3_stage_124 <= bright_bright_update_0_write_write_3_stage_123;
      bright_bright_update_0_write_write_3_stage_125 <= bright_bright_update_0_write_write_3_stage_124;
      bright_bright_update_0_write_write_3_stage_126 <= bright_bright_update_0_write_write_3_stage_125;
      bright_bright_update_0_write_write_3_stage_127 <= bright_bright_update_0_write_write_3_stage_126;
      bright_bright_update_0_write_write_3_stage_128 <= bright_bright_update_0_write_write_3_stage_127;
      bright_bright_update_0_write_write_3_stage_129 <= bright_bright_update_0_write_write_3_stage_128;
      bright_bright_update_0_write_write_3_stage_130 <= bright_bright_update_0_write_write_3_stage_129;
      bright_bright_update_0_write_write_3_stage_131 <= bright_bright_update_0_write_write_3_stage_130;
      bright_bright_update_0_write_write_3_stage_132 <= bright_bright_update_0_write_write_3_stage_131;
      bright_bright_update_0_write_write_3_stage_133 <= bright_bright_update_0_write_write_3_stage_132;
      bright_bright_update_0_write_write_3_stage_134 <= bright_bright_update_0_write_write_3_stage_133;
      bright_bright_update_0_write_write_3_stage_135 <= bright_bright_update_0_write_write_3_stage_134;
      bright_bright_update_0_write_write_3_stage_136 <= bright_bright_update_0_write_write_3_stage_135;
      bright_bright_update_0_write_write_3_stage_137 <= bright_bright_update_0_write_write_3_stage_136;
      bright_bright_update_0_write_write_3_stage_138 <= bright_bright_update_0_write_write_3_stage_137;
      bright_bright_update_0_write_write_3_stage_139 <= bright_bright_update_0_write_write_3_stage_138;
      bright_bright_update_0_write_write_3_stage_140 <= bright_bright_update_0_write_write_3_stage_139;
      bright_bright_update_0_write_write_3_stage_141 <= bright_bright_update_0_write_write_3_stage_140;
      bright_bright_update_0_write_write_3_stage_142 <= bright_bright_update_0_write_write_3_stage_141;
      bright_bright_update_0_write_write_3_stage_143 <= bright_bright_update_0_write_write_3_stage_142;
      bright_bright_update_0_write_write_3_stage_144 <= bright_bright_update_0_write_write_3_stage_143;
      bright_bright_update_0_write_write_3_stage_145 <= bright_bright_update_0_write_write_3_stage_144;
      bright_bright_update_0_write_write_3_stage_146 <= bright_bright_update_0_write_write_3_stage_145;
      bright_bright_update_0_write_write_3_stage_147 <= bright_bright_update_0_write_write_3_stage_146;
      bright_bright_update_0_write_write_3_stage_148 <= bright_bright_update_0_write_write_3_stage_147;
      bright_bright_update_0_write_write_3_stage_149 <= bright_bright_update_0_write_write_3_stage_148;
      bright_bright_update_0_write_write_3_stage_150 <= bright_bright_update_0_write_write_3_stage_149;
      bright_bright_update_0_write_write_3_stage_151 <= bright_bright_update_0_write_write_3_stage_150;
      bright_bright_update_0_write_write_3_stage_152 <= bright_bright_update_0_write_write_3_stage_151;
      bright_bright_update_0_write_write_3_stage_153 <= bright_bright_update_0_write_write_3_stage_152;
      bright_bright_update_0_write_write_3_stage_154 <= bright_bright_update_0_write_write_3_stage_153;
      bright_bright_update_0_write_write_3_stage_155 <= bright_bright_update_0_write_write_3_stage_154;
      bright_bright_update_0_write_write_3_stage_156 <= bright_bright_update_0_write_write_3_stage_155;
      bright_bright_update_0_write_write_3_stage_157 <= bright_bright_update_0_write_write_3_stage_156;
      bright_bright_update_0_write_write_3_stage_158 <= bright_bright_update_0_write_write_3_stage_157;
      bright_bright_update_0_write_write_3_stage_159 <= bright_bright_update_0_write_write_3_stage_158;
      bright_bright_update_0_write_write_3_stage_160 <= bright_bright_update_0_write_write_3_stage_159;
      bright_bright_update_0_write_write_3_stage_161 <= bright_bright_update_0_write_write_3_stage_160;
      bright_bright_update_0_write_write_3_stage_162 <= bright_bright_update_0_write_write_3_stage_161;
      bright_bright_update_0_write_write_3_stage_163 <= bright_bright_update_0_write_write_3_stage_162;
      bright_bright_update_0_write_write_3_stage_164 <= bright_bright_update_0_write_write_3_stage_163;
      bright_bright_update_0_write_write_3_stage_165 <= bright_bright_update_0_write_write_3_stage_164;
      bright_bright_update_0_write_write_3_stage_166 <= bright_bright_update_0_write_write_3_stage_165;
      bright_bright_update_0_write_write_3_stage_167 <= bright_bright_update_0_write_write_3_stage_166;
      bright_bright_update_0_write_write_3_stage_168 <= bright_bright_update_0_write_write_3_stage_167;
      bright_bright_update_0_write_write_3_stage_169 <= bright_bright_update_0_write_write_3_stage_168;
      bright_bright_update_0_write_write_3_stage_170 <= bright_bright_update_0_write_write_3_stage_169;
      bright_bright_update_0_write_write_3_stage_171 <= bright_bright_update_0_write_write_3_stage_170;
      bright_bright_update_0_write_write_3_stage_172 <= bright_bright_update_0_write_write_3_stage_171;
      bright_bright_update_0_write_write_3_stage_173 <= bright_bright_update_0_write_write_3_stage_172;
      bright_bright_update_0_write_write_3_stage_174 <= bright_bright_update_0_write_write_3_stage_173;
      bright_bright_update_0_write_write_3_stage_175 <= bright_bright_update_0_write_write_3_stage_174;
      bright_bright_update_0_write_write_3_stage_176 <= bright_bright_update_0_write_write_3_stage_175;
      bright_bright_update_0_write_write_3_stage_177 <= bright_bright_update_0_write_write_3_stage_176;
      bright_bright_update_0_write_write_3_stage_178 <= bright_bright_update_0_write_write_3_stage_177;
      bright_bright_update_0_write_write_3_stage_179 <= bright_bright_update_0_write_write_3_stage_178;
      bright_bright_update_0_write_write_3_stage_180 <= bright_bright_update_0_write_write_3_stage_179;
      bright_bright_update_0_write_write_3_stage_181 <= bright_bright_update_0_write_write_3_stage_180;
      in_dark_update_0_read_read_6_stage_11 <= in_dark_update_0_read_read_6;
      in_dark_update_0_read_read_6_stage_12 <= in_dark_update_0_read_read_6_stage_11;
      in_dark_update_0_read_read_6_stage_13 <= in_dark_update_0_read_read_6_stage_12;
      in_dark_update_0_read_read_6_stage_14 <= in_dark_update_0_read_read_6_stage_13;
      in_dark_update_0_read_read_6_stage_15 <= in_dark_update_0_read_read_6_stage_14;
      in_dark_update_0_read_read_6_stage_16 <= in_dark_update_0_read_read_6_stage_15;
      in_dark_update_0_read_read_6_stage_17 <= in_dark_update_0_read_read_6_stage_16;
      in_dark_update_0_read_read_6_stage_18 <= in_dark_update_0_read_read_6_stage_17;
      in_dark_update_0_read_read_6_stage_19 <= in_dark_update_0_read_read_6_stage_18;
      in_dark_update_0_read_read_6_stage_20 <= in_dark_update_0_read_read_6_stage_19;
      in_dark_update_0_read_read_6_stage_21 <= in_dark_update_0_read_read_6_stage_20;
      in_dark_update_0_read_read_6_stage_22 <= in_dark_update_0_read_read_6_stage_21;
      in_dark_update_0_read_read_6_stage_23 <= in_dark_update_0_read_read_6_stage_22;
      in_dark_update_0_read_read_6_stage_24 <= in_dark_update_0_read_read_6_stage_23;
      in_dark_update_0_read_read_6_stage_25 <= in_dark_update_0_read_read_6_stage_24;
      in_dark_update_0_read_read_6_stage_26 <= in_dark_update_0_read_read_6_stage_25;
      in_dark_update_0_read_read_6_stage_27 <= in_dark_update_0_read_read_6_stage_26;
      in_dark_update_0_read_read_6_stage_28 <= in_dark_update_0_read_read_6_stage_27;
      in_dark_update_0_read_read_6_stage_29 <= in_dark_update_0_read_read_6_stage_28;
      in_dark_update_0_read_read_6_stage_30 <= in_dark_update_0_read_read_6_stage_29;
      in_dark_update_0_read_read_6_stage_31 <= in_dark_update_0_read_read_6_stage_30;
      in_dark_update_0_read_read_6_stage_32 <= in_dark_update_0_read_read_6_stage_31;
      in_dark_update_0_read_read_6_stage_33 <= in_dark_update_0_read_read_6_stage_32;
      in_dark_update_0_read_read_6_stage_34 <= in_dark_update_0_read_read_6_stage_33;
      in_dark_update_0_read_read_6_stage_35 <= in_dark_update_0_read_read_6_stage_34;
      in_dark_update_0_read_read_6_stage_36 <= in_dark_update_0_read_read_6_stage_35;
      in_dark_update_0_read_read_6_stage_37 <= in_dark_update_0_read_read_6_stage_36;
      in_dark_update_0_read_read_6_stage_38 <= in_dark_update_0_read_read_6_stage_37;
      in_dark_update_0_read_read_6_stage_39 <= in_dark_update_0_read_read_6_stage_38;
      in_dark_update_0_read_read_6_stage_40 <= in_dark_update_0_read_read_6_stage_39;
      in_dark_update_0_read_read_6_stage_41 <= in_dark_update_0_read_read_6_stage_40;
      in_dark_update_0_read_read_6_stage_42 <= in_dark_update_0_read_read_6_stage_41;
      in_dark_update_0_read_read_6_stage_43 <= in_dark_update_0_read_read_6_stage_42;
      in_dark_update_0_read_read_6_stage_44 <= in_dark_update_0_read_read_6_stage_43;
      in_dark_update_0_read_read_6_stage_45 <= in_dark_update_0_read_read_6_stage_44;
      in_dark_update_0_read_read_6_stage_46 <= in_dark_update_0_read_read_6_stage_45;
      in_dark_update_0_read_read_6_stage_47 <= in_dark_update_0_read_read_6_stage_46;
      in_dark_update_0_read_read_6_stage_48 <= in_dark_update_0_read_read_6_stage_47;
      in_dark_update_0_read_read_6_stage_49 <= in_dark_update_0_read_read_6_stage_48;
      in_dark_update_0_read_read_6_stage_50 <= in_dark_update_0_read_read_6_stage_49;
      in_dark_update_0_read_read_6_stage_51 <= in_dark_update_0_read_read_6_stage_50;
      in_dark_update_0_read_read_6_stage_52 <= in_dark_update_0_read_read_6_stage_51;
      in_dark_update_0_read_read_6_stage_53 <= in_dark_update_0_read_read_6_stage_52;
      in_dark_update_0_read_read_6_stage_54 <= in_dark_update_0_read_read_6_stage_53;
      in_dark_update_0_read_read_6_stage_55 <= in_dark_update_0_read_read_6_stage_54;
      in_dark_update_0_read_read_6_stage_56 <= in_dark_update_0_read_read_6_stage_55;
      in_dark_update_0_read_read_6_stage_57 <= in_dark_update_0_read_read_6_stage_56;
      in_dark_update_0_read_read_6_stage_58 <= in_dark_update_0_read_read_6_stage_57;
      in_dark_update_0_read_read_6_stage_59 <= in_dark_update_0_read_read_6_stage_58;
      in_dark_update_0_read_read_6_stage_60 <= in_dark_update_0_read_read_6_stage_59;
      in_dark_update_0_read_read_6_stage_61 <= in_dark_update_0_read_read_6_stage_60;
      in_dark_update_0_read_read_6_stage_62 <= in_dark_update_0_read_read_6_stage_61;
      in_dark_update_0_read_read_6_stage_63 <= in_dark_update_0_read_read_6_stage_62;
      in_dark_update_0_read_read_6_stage_64 <= in_dark_update_0_read_read_6_stage_63;
      in_dark_update_0_read_read_6_stage_65 <= in_dark_update_0_read_read_6_stage_64;
      in_dark_update_0_read_read_6_stage_66 <= in_dark_update_0_read_read_6_stage_65;
      in_dark_update_0_read_read_6_stage_67 <= in_dark_update_0_read_read_6_stage_66;
      in_dark_update_0_read_read_6_stage_68 <= in_dark_update_0_read_read_6_stage_67;
      in_dark_update_0_read_read_6_stage_69 <= in_dark_update_0_read_read_6_stage_68;
      in_dark_update_0_read_read_6_stage_70 <= in_dark_update_0_read_read_6_stage_69;
      in_dark_update_0_read_read_6_stage_71 <= in_dark_update_0_read_read_6_stage_70;
      in_dark_update_0_read_read_6_stage_72 <= in_dark_update_0_read_read_6_stage_71;
      in_dark_update_0_read_read_6_stage_73 <= in_dark_update_0_read_read_6_stage_72;
      in_dark_update_0_read_read_6_stage_74 <= in_dark_update_0_read_read_6_stage_73;
      in_dark_update_0_read_read_6_stage_75 <= in_dark_update_0_read_read_6_stage_74;
      in_dark_update_0_read_read_6_stage_76 <= in_dark_update_0_read_read_6_stage_75;
      in_dark_update_0_read_read_6_stage_77 <= in_dark_update_0_read_read_6_stage_76;
      in_dark_update_0_read_read_6_stage_78 <= in_dark_update_0_read_read_6_stage_77;
      in_dark_update_0_read_read_6_stage_79 <= in_dark_update_0_read_read_6_stage_78;
      in_dark_update_0_read_read_6_stage_80 <= in_dark_update_0_read_read_6_stage_79;
      in_dark_update_0_read_read_6_stage_81 <= in_dark_update_0_read_read_6_stage_80;
      in_dark_update_0_read_read_6_stage_82 <= in_dark_update_0_read_read_6_stage_81;
      in_dark_update_0_read_read_6_stage_83 <= in_dark_update_0_read_read_6_stage_82;
      in_dark_update_0_read_read_6_stage_84 <= in_dark_update_0_read_read_6_stage_83;
      in_dark_update_0_read_read_6_stage_85 <= in_dark_update_0_read_read_6_stage_84;
      in_dark_update_0_read_read_6_stage_86 <= in_dark_update_0_read_read_6_stage_85;
      in_dark_update_0_read_read_6_stage_87 <= in_dark_update_0_read_read_6_stage_86;
      in_dark_update_0_read_read_6_stage_88 <= in_dark_update_0_read_read_6_stage_87;
      in_dark_update_0_read_read_6_stage_89 <= in_dark_update_0_read_read_6_stage_88;
      in_dark_update_0_read_read_6_stage_90 <= in_dark_update_0_read_read_6_stage_89;
      in_dark_update_0_read_read_6_stage_91 <= in_dark_update_0_read_read_6_stage_90;
      in_dark_update_0_read_read_6_stage_92 <= in_dark_update_0_read_read_6_stage_91;
      in_dark_update_0_read_read_6_stage_93 <= in_dark_update_0_read_read_6_stage_92;
      in_dark_update_0_read_read_6_stage_94 <= in_dark_update_0_read_read_6_stage_93;
      in_dark_update_0_read_read_6_stage_95 <= in_dark_update_0_read_read_6_stage_94;
      in_dark_update_0_read_read_6_stage_96 <= in_dark_update_0_read_read_6_stage_95;
      in_dark_update_0_read_read_6_stage_97 <= in_dark_update_0_read_read_6_stage_96;
      in_dark_update_0_read_read_6_stage_98 <= in_dark_update_0_read_read_6_stage_97;
      in_dark_update_0_read_read_6_stage_99 <= in_dark_update_0_read_read_6_stage_98;
      in_dark_update_0_read_read_6_stage_100 <= in_dark_update_0_read_read_6_stage_99;
      in_dark_update_0_read_read_6_stage_101 <= in_dark_update_0_read_read_6_stage_100;
      in_dark_update_0_read_read_6_stage_102 <= in_dark_update_0_read_read_6_stage_101;
      in_dark_update_0_read_read_6_stage_103 <= in_dark_update_0_read_read_6_stage_102;
      in_dark_update_0_read_read_6_stage_104 <= in_dark_update_0_read_read_6_stage_103;
      in_dark_update_0_read_read_6_stage_105 <= in_dark_update_0_read_read_6_stage_104;
      in_dark_update_0_read_read_6_stage_106 <= in_dark_update_0_read_read_6_stage_105;
      in_dark_update_0_read_read_6_stage_107 <= in_dark_update_0_read_read_6_stage_106;
      in_dark_update_0_read_read_6_stage_108 <= in_dark_update_0_read_read_6_stage_107;
      in_dark_update_0_read_read_6_stage_109 <= in_dark_update_0_read_read_6_stage_108;
      in_dark_update_0_read_read_6_stage_110 <= in_dark_update_0_read_read_6_stage_109;
      in_dark_update_0_read_read_6_stage_111 <= in_dark_update_0_read_read_6_stage_110;
      in_dark_update_0_read_read_6_stage_112 <= in_dark_update_0_read_read_6_stage_111;
      in_dark_update_0_read_read_6_stage_113 <= in_dark_update_0_read_read_6_stage_112;
      in_dark_update_0_read_read_6_stage_114 <= in_dark_update_0_read_read_6_stage_113;
      in_dark_update_0_read_read_6_stage_115 <= in_dark_update_0_read_read_6_stage_114;
      in_dark_update_0_read_read_6_stage_116 <= in_dark_update_0_read_read_6_stage_115;
      in_dark_update_0_read_read_6_stage_117 <= in_dark_update_0_read_read_6_stage_116;
      in_dark_update_0_read_read_6_stage_118 <= in_dark_update_0_read_read_6_stage_117;
      in_dark_update_0_read_read_6_stage_119 <= in_dark_update_0_read_read_6_stage_118;
      in_dark_update_0_read_read_6_stage_120 <= in_dark_update_0_read_read_6_stage_119;
      in_dark_update_0_read_read_6_stage_121 <= in_dark_update_0_read_read_6_stage_120;
      in_dark_update_0_read_read_6_stage_122 <= in_dark_update_0_read_read_6_stage_121;
      in_dark_update_0_read_read_6_stage_123 <= in_dark_update_0_read_read_6_stage_122;
      in_dark_update_0_read_read_6_stage_124 <= in_dark_update_0_read_read_6_stage_123;
      in_dark_update_0_read_read_6_stage_125 <= in_dark_update_0_read_read_6_stage_124;
      in_dark_update_0_read_read_6_stage_126 <= in_dark_update_0_read_read_6_stage_125;
      in_dark_update_0_read_read_6_stage_127 <= in_dark_update_0_read_read_6_stage_126;
      in_dark_update_0_read_read_6_stage_128 <= in_dark_update_0_read_read_6_stage_127;
      in_dark_update_0_read_read_6_stage_129 <= in_dark_update_0_read_read_6_stage_128;
      in_dark_update_0_read_read_6_stage_130 <= in_dark_update_0_read_read_6_stage_129;
      in_dark_update_0_read_read_6_stage_131 <= in_dark_update_0_read_read_6_stage_130;
      in_dark_update_0_read_read_6_stage_132 <= in_dark_update_0_read_read_6_stage_131;
      in_dark_update_0_read_read_6_stage_133 <= in_dark_update_0_read_read_6_stage_132;
      in_dark_update_0_read_read_6_stage_134 <= in_dark_update_0_read_read_6_stage_133;
      in_dark_update_0_read_read_6_stage_135 <= in_dark_update_0_read_read_6_stage_134;
      in_dark_update_0_read_read_6_stage_136 <= in_dark_update_0_read_read_6_stage_135;
      in_dark_update_0_read_read_6_stage_137 <= in_dark_update_0_read_read_6_stage_136;
      in_dark_update_0_read_read_6_stage_138 <= in_dark_update_0_read_read_6_stage_137;
      in_dark_update_0_read_read_6_stage_139 <= in_dark_update_0_read_read_6_stage_138;
      in_dark_update_0_read_read_6_stage_140 <= in_dark_update_0_read_read_6_stage_139;
      in_dark_update_0_read_read_6_stage_141 <= in_dark_update_0_read_read_6_stage_140;
      in_dark_update_0_read_read_6_stage_142 <= in_dark_update_0_read_read_6_stage_141;
      in_dark_update_0_read_read_6_stage_143 <= in_dark_update_0_read_read_6_stage_142;
      in_dark_update_0_read_read_6_stage_144 <= in_dark_update_0_read_read_6_stage_143;
      in_dark_update_0_read_read_6_stage_145 <= in_dark_update_0_read_read_6_stage_144;
      in_dark_update_0_read_read_6_stage_146 <= in_dark_update_0_read_read_6_stage_145;
      in_dark_update_0_read_read_6_stage_147 <= in_dark_update_0_read_read_6_stage_146;
      in_dark_update_0_read_read_6_stage_148 <= in_dark_update_0_read_read_6_stage_147;
      in_dark_update_0_read_read_6_stage_149 <= in_dark_update_0_read_read_6_stage_148;
      in_dark_update_0_read_read_6_stage_150 <= in_dark_update_0_read_read_6_stage_149;
      in_dark_update_0_read_read_6_stage_151 <= in_dark_update_0_read_read_6_stage_150;
      in_dark_update_0_read_read_6_stage_152 <= in_dark_update_0_read_read_6_stage_151;
      in_dark_update_0_read_read_6_stage_153 <= in_dark_update_0_read_read_6_stage_152;
      in_dark_update_0_read_read_6_stage_154 <= in_dark_update_0_read_read_6_stage_153;
      in_dark_update_0_read_read_6_stage_155 <= in_dark_update_0_read_read_6_stage_154;
      in_dark_update_0_read_read_6_stage_156 <= in_dark_update_0_read_read_6_stage_155;
      in_dark_update_0_read_read_6_stage_157 <= in_dark_update_0_read_read_6_stage_156;
      in_dark_update_0_read_read_6_stage_158 <= in_dark_update_0_read_read_6_stage_157;
      in_dark_update_0_read_read_6_stage_159 <= in_dark_update_0_read_read_6_stage_158;
      in_dark_update_0_read_read_6_stage_160 <= in_dark_update_0_read_read_6_stage_159;
      in_dark_update_0_read_read_6_stage_161 <= in_dark_update_0_read_read_6_stage_160;
      in_dark_update_0_read_read_6_stage_162 <= in_dark_update_0_read_read_6_stage_161;
      in_dark_update_0_read_read_6_stage_163 <= in_dark_update_0_read_read_6_stage_162;
      in_dark_update_0_read_read_6_stage_164 <= in_dark_update_0_read_read_6_stage_163;
      in_dark_update_0_read_read_6_stage_165 <= in_dark_update_0_read_read_6_stage_164;
      in_dark_update_0_read_read_6_stage_166 <= in_dark_update_0_read_read_6_stage_165;
      in_dark_update_0_read_read_6_stage_167 <= in_dark_update_0_read_read_6_stage_166;
      in_dark_update_0_read_read_6_stage_168 <= in_dark_update_0_read_read_6_stage_167;
      in_dark_update_0_read_read_6_stage_169 <= in_dark_update_0_read_read_6_stage_168;
      in_dark_update_0_read_read_6_stage_170 <= in_dark_update_0_read_read_6_stage_169;
      in_dark_update_0_read_read_6_stage_171 <= in_dark_update_0_read_read_6_stage_170;
      in_dark_update_0_read_read_6_stage_172 <= in_dark_update_0_read_read_6_stage_171;
      in_dark_update_0_read_read_6_stage_173 <= in_dark_update_0_read_read_6_stage_172;
      in_dark_update_0_read_read_6_stage_174 <= in_dark_update_0_read_read_6_stage_173;
      in_dark_update_0_read_read_6_stage_175 <= in_dark_update_0_read_read_6_stage_174;
      in_dark_update_0_read_read_6_stage_176 <= in_dark_update_0_read_read_6_stage_175;
      in_dark_update_0_read_read_6_stage_177 <= in_dark_update_0_read_read_6_stage_176;
      in_dark_update_0_read_read_6_stage_178 <= in_dark_update_0_read_read_6_stage_177;
      in_dark_update_0_read_read_6_stage_179 <= in_dark_update_0_read_read_6_stage_178;
      in_dark_update_0_read_read_6_stage_180 <= in_dark_update_0_read_read_6_stage_179;
      in_dark_update_0_read_read_6_stage_181 <= in_dark_update_0_read_read_6_stage_180;
      dark_update_0_stage_12 <= dark_update_0;
      dark_update_0_stage_13 <= dark_update_0_stage_12;
      dark_update_0_stage_14 <= dark_update_0_stage_13;
      dark_update_0_stage_15 <= dark_update_0_stage_14;
      dark_update_0_stage_16 <= dark_update_0_stage_15;
      dark_update_0_stage_17 <= dark_update_0_stage_16;
      dark_update_0_stage_18 <= dark_update_0_stage_17;
      dark_update_0_stage_19 <= dark_update_0_stage_18;
      dark_update_0_stage_20 <= dark_update_0_stage_19;
      dark_update_0_stage_21 <= dark_update_0_stage_20;
      dark_update_0_stage_22 <= dark_update_0_stage_21;
      dark_update_0_stage_23 <= dark_update_0_stage_22;
      dark_update_0_stage_24 <= dark_update_0_stage_23;
      dark_update_0_stage_25 <= dark_update_0_stage_24;
      dark_update_0_stage_26 <= dark_update_0_stage_25;
      dark_update_0_stage_27 <= dark_update_0_stage_26;
      dark_update_0_stage_28 <= dark_update_0_stage_27;
      dark_update_0_stage_29 <= dark_update_0_stage_28;
      dark_update_0_stage_30 <= dark_update_0_stage_29;
      dark_update_0_stage_31 <= dark_update_0_stage_30;
      dark_update_0_stage_32 <= dark_update_0_stage_31;
      dark_update_0_stage_33 <= dark_update_0_stage_32;
      dark_update_0_stage_34 <= dark_update_0_stage_33;
      dark_update_0_stage_35 <= dark_update_0_stage_34;
      dark_update_0_stage_36 <= dark_update_0_stage_35;
      dark_update_0_stage_37 <= dark_update_0_stage_36;
      dark_update_0_stage_38 <= dark_update_0_stage_37;
      dark_update_0_stage_39 <= dark_update_0_stage_38;
      dark_update_0_stage_40 <= dark_update_0_stage_39;
      dark_update_0_stage_41 <= dark_update_0_stage_40;
      dark_update_0_stage_42 <= dark_update_0_stage_41;
      dark_update_0_stage_43 <= dark_update_0_stage_42;
      dark_update_0_stage_44 <= dark_update_0_stage_43;
      dark_update_0_stage_45 <= dark_update_0_stage_44;
      dark_update_0_stage_46 <= dark_update_0_stage_45;
      dark_update_0_stage_47 <= dark_update_0_stage_46;
      dark_update_0_stage_48 <= dark_update_0_stage_47;
      dark_update_0_stage_49 <= dark_update_0_stage_48;
      dark_update_0_stage_50 <= dark_update_0_stage_49;
      dark_update_0_stage_51 <= dark_update_0_stage_50;
      dark_update_0_stage_52 <= dark_update_0_stage_51;
      dark_update_0_stage_53 <= dark_update_0_stage_52;
      dark_update_0_stage_54 <= dark_update_0_stage_53;
      dark_update_0_stage_55 <= dark_update_0_stage_54;
      dark_update_0_stage_56 <= dark_update_0_stage_55;
      dark_update_0_stage_57 <= dark_update_0_stage_56;
      dark_update_0_stage_58 <= dark_update_0_stage_57;
      dark_update_0_stage_59 <= dark_update_0_stage_58;
      dark_update_0_stage_60 <= dark_update_0_stage_59;
      dark_update_0_stage_61 <= dark_update_0_stage_60;
      dark_update_0_stage_62 <= dark_update_0_stage_61;
      dark_update_0_stage_63 <= dark_update_0_stage_62;
      dark_update_0_stage_64 <= dark_update_0_stage_63;
      dark_update_0_stage_65 <= dark_update_0_stage_64;
      dark_update_0_stage_66 <= dark_update_0_stage_65;
      dark_update_0_stage_67 <= dark_update_0_stage_66;
      dark_update_0_stage_68 <= dark_update_0_stage_67;
      dark_update_0_stage_69 <= dark_update_0_stage_68;
      dark_update_0_stage_70 <= dark_update_0_stage_69;
      dark_update_0_stage_71 <= dark_update_0_stage_70;
      dark_update_0_stage_72 <= dark_update_0_stage_71;
      dark_update_0_stage_73 <= dark_update_0_stage_72;
      dark_update_0_stage_74 <= dark_update_0_stage_73;
      dark_update_0_stage_75 <= dark_update_0_stage_74;
      dark_update_0_stage_76 <= dark_update_0_stage_75;
      dark_update_0_stage_77 <= dark_update_0_stage_76;
      dark_update_0_stage_78 <= dark_update_0_stage_77;
      dark_update_0_stage_79 <= dark_update_0_stage_78;
      dark_update_0_stage_80 <= dark_update_0_stage_79;
      dark_update_0_stage_81 <= dark_update_0_stage_80;
      dark_update_0_stage_82 <= dark_update_0_stage_81;
      dark_update_0_stage_83 <= dark_update_0_stage_82;
      dark_update_0_stage_84 <= dark_update_0_stage_83;
      dark_update_0_stage_85 <= dark_update_0_stage_84;
      dark_update_0_stage_86 <= dark_update_0_stage_85;
      dark_update_0_stage_87 <= dark_update_0_stage_86;
      dark_update_0_stage_88 <= dark_update_0_stage_87;
      dark_update_0_stage_89 <= dark_update_0_stage_88;
      dark_update_0_stage_90 <= dark_update_0_stage_89;
      dark_update_0_stage_91 <= dark_update_0_stage_90;
      dark_update_0_stage_92 <= dark_update_0_stage_91;
      dark_update_0_stage_93 <= dark_update_0_stage_92;
      dark_update_0_stage_94 <= dark_update_0_stage_93;
      dark_update_0_stage_95 <= dark_update_0_stage_94;
      dark_update_0_stage_96 <= dark_update_0_stage_95;
      dark_update_0_stage_97 <= dark_update_0_stage_96;
      dark_update_0_stage_98 <= dark_update_0_stage_97;
      dark_update_0_stage_99 <= dark_update_0_stage_98;
      dark_update_0_stage_100 <= dark_update_0_stage_99;
      dark_update_0_stage_101 <= dark_update_0_stage_100;
      dark_update_0_stage_102 <= dark_update_0_stage_101;
      dark_update_0_stage_103 <= dark_update_0_stage_102;
      dark_update_0_stage_104 <= dark_update_0_stage_103;
      dark_update_0_stage_105 <= dark_update_0_stage_104;
      dark_update_0_stage_106 <= dark_update_0_stage_105;
      dark_update_0_stage_107 <= dark_update_0_stage_106;
      dark_update_0_stage_108 <= dark_update_0_stage_107;
      dark_update_0_stage_109 <= dark_update_0_stage_108;
      dark_update_0_stage_110 <= dark_update_0_stage_109;
      dark_update_0_stage_111 <= dark_update_0_stage_110;
      dark_update_0_stage_112 <= dark_update_0_stage_111;
      dark_update_0_stage_113 <= dark_update_0_stage_112;
      dark_update_0_stage_114 <= dark_update_0_stage_113;
      dark_update_0_stage_115 <= dark_update_0_stage_114;
      dark_update_0_stage_116 <= dark_update_0_stage_115;
      dark_update_0_stage_117 <= dark_update_0_stage_116;
      dark_update_0_stage_118 <= dark_update_0_stage_117;
      dark_update_0_stage_119 <= dark_update_0_stage_118;
      dark_update_0_stage_120 <= dark_update_0_stage_119;
      dark_update_0_stage_121 <= dark_update_0_stage_120;
      dark_update_0_stage_122 <= dark_update_0_stage_121;
      dark_update_0_stage_123 <= dark_update_0_stage_122;
      dark_update_0_stage_124 <= dark_update_0_stage_123;
      dark_update_0_stage_125 <= dark_update_0_stage_124;
      dark_update_0_stage_126 <= dark_update_0_stage_125;
      dark_update_0_stage_127 <= dark_update_0_stage_126;
      dark_update_0_stage_128 <= dark_update_0_stage_127;
      dark_update_0_stage_129 <= dark_update_0_stage_128;
      dark_update_0_stage_130 <= dark_update_0_stage_129;
      dark_update_0_stage_131 <= dark_update_0_stage_130;
      dark_update_0_stage_132 <= dark_update_0_stage_131;
      dark_update_0_stage_133 <= dark_update_0_stage_132;
      dark_update_0_stage_134 <= dark_update_0_stage_133;
      dark_update_0_stage_135 <= dark_update_0_stage_134;
      dark_update_0_stage_136 <= dark_update_0_stage_135;
      dark_update_0_stage_137 <= dark_update_0_stage_136;
      dark_update_0_stage_138 <= dark_update_0_stage_137;
      dark_update_0_stage_139 <= dark_update_0_stage_138;
      dark_update_0_stage_140 <= dark_update_0_stage_139;
      dark_update_0_stage_141 <= dark_update_0_stage_140;
      dark_update_0_stage_142 <= dark_update_0_stage_141;
      dark_update_0_stage_143 <= dark_update_0_stage_142;
      dark_update_0_stage_144 <= dark_update_0_stage_143;
      dark_update_0_stage_145 <= dark_update_0_stage_144;
      dark_update_0_stage_146 <= dark_update_0_stage_145;
      dark_update_0_stage_147 <= dark_update_0_stage_146;
      dark_update_0_stage_148 <= dark_update_0_stage_147;
      dark_update_0_stage_149 <= dark_update_0_stage_148;
      dark_update_0_stage_150 <= dark_update_0_stage_149;
      dark_update_0_stage_151 <= dark_update_0_stage_150;
      dark_update_0_stage_152 <= dark_update_0_stage_151;
      dark_update_0_stage_153 <= dark_update_0_stage_152;
      dark_update_0_stage_154 <= dark_update_0_stage_153;
      dark_update_0_stage_155 <= dark_update_0_stage_154;
      dark_update_0_stage_156 <= dark_update_0_stage_155;
      dark_update_0_stage_157 <= dark_update_0_stage_156;
      dark_update_0_stage_158 <= dark_update_0_stage_157;
      dark_update_0_stage_159 <= dark_update_0_stage_158;
      dark_update_0_stage_160 <= dark_update_0_stage_159;
      dark_update_0_stage_161 <= dark_update_0_stage_160;
      dark_update_0_stage_162 <= dark_update_0_stage_161;
      dark_update_0_stage_163 <= dark_update_0_stage_162;
      dark_update_0_stage_164 <= dark_update_0_stage_163;
      dark_update_0_stage_165 <= dark_update_0_stage_164;
      dark_update_0_stage_166 <= dark_update_0_stage_165;
      dark_update_0_stage_167 <= dark_update_0_stage_166;
      dark_update_0_stage_168 <= dark_update_0_stage_167;
      dark_update_0_stage_169 <= dark_update_0_stage_168;
      dark_update_0_stage_170 <= dark_update_0_stage_169;
      dark_update_0_stage_171 <= dark_update_0_stage_170;
      dark_update_0_stage_172 <= dark_update_0_stage_171;
      dark_update_0_stage_173 <= dark_update_0_stage_172;
      dark_update_0_stage_174 <= dark_update_0_stage_173;
      dark_update_0_stage_175 <= dark_update_0_stage_174;
      dark_update_0_stage_176 <= dark_update_0_stage_175;
      dark_update_0_stage_177 <= dark_update_0_stage_176;
      dark_update_0_stage_178 <= dark_update_0_stage_177;
      dark_update_0_stage_179 <= dark_update_0_stage_178;
      dark_update_0_stage_180 <= dark_update_0_stage_179;
      dark_update_0_stage_181 <= dark_update_0_stage_180;
      dark_dark_update_0_write_write_7_stage_13 <= dark_dark_update_0_write_write_7;
      dark_dark_update_0_write_write_7_stage_14 <= dark_dark_update_0_write_write_7_stage_13;
      dark_dark_update_0_write_write_7_stage_15 <= dark_dark_update_0_write_write_7_stage_14;
      dark_dark_update_0_write_write_7_stage_16 <= dark_dark_update_0_write_write_7_stage_15;
      dark_dark_update_0_write_write_7_stage_17 <= dark_dark_update_0_write_write_7_stage_16;
      dark_dark_update_0_write_write_7_stage_18 <= dark_dark_update_0_write_write_7_stage_17;
      dark_dark_update_0_write_write_7_stage_19 <= dark_dark_update_0_write_write_7_stage_18;
      dark_dark_update_0_write_write_7_stage_20 <= dark_dark_update_0_write_write_7_stage_19;
      dark_dark_update_0_write_write_7_stage_21 <= dark_dark_update_0_write_write_7_stage_20;
      dark_dark_update_0_write_write_7_stage_22 <= dark_dark_update_0_write_write_7_stage_21;
      dark_dark_update_0_write_write_7_stage_23 <= dark_dark_update_0_write_write_7_stage_22;
      dark_dark_update_0_write_write_7_stage_24 <= dark_dark_update_0_write_write_7_stage_23;
      dark_dark_update_0_write_write_7_stage_25 <= dark_dark_update_0_write_write_7_stage_24;
      dark_dark_update_0_write_write_7_stage_26 <= dark_dark_update_0_write_write_7_stage_25;
      dark_dark_update_0_write_write_7_stage_27 <= dark_dark_update_0_write_write_7_stage_26;
      dark_dark_update_0_write_write_7_stage_28 <= dark_dark_update_0_write_write_7_stage_27;
      dark_dark_update_0_write_write_7_stage_29 <= dark_dark_update_0_write_write_7_stage_28;
      dark_dark_update_0_write_write_7_stage_30 <= dark_dark_update_0_write_write_7_stage_29;
      dark_dark_update_0_write_write_7_stage_31 <= dark_dark_update_0_write_write_7_stage_30;
      dark_dark_update_0_write_write_7_stage_32 <= dark_dark_update_0_write_write_7_stage_31;
      dark_dark_update_0_write_write_7_stage_33 <= dark_dark_update_0_write_write_7_stage_32;
      dark_dark_update_0_write_write_7_stage_34 <= dark_dark_update_0_write_write_7_stage_33;
      dark_dark_update_0_write_write_7_stage_35 <= dark_dark_update_0_write_write_7_stage_34;
      dark_dark_update_0_write_write_7_stage_36 <= dark_dark_update_0_write_write_7_stage_35;
      dark_dark_update_0_write_write_7_stage_37 <= dark_dark_update_0_write_write_7_stage_36;
      dark_dark_update_0_write_write_7_stage_38 <= dark_dark_update_0_write_write_7_stage_37;
      dark_dark_update_0_write_write_7_stage_39 <= dark_dark_update_0_write_write_7_stage_38;
      dark_dark_update_0_write_write_7_stage_40 <= dark_dark_update_0_write_write_7_stage_39;
      dark_dark_update_0_write_write_7_stage_41 <= dark_dark_update_0_write_write_7_stage_40;
      dark_dark_update_0_write_write_7_stage_42 <= dark_dark_update_0_write_write_7_stage_41;
      dark_dark_update_0_write_write_7_stage_43 <= dark_dark_update_0_write_write_7_stage_42;
      dark_dark_update_0_write_write_7_stage_44 <= dark_dark_update_0_write_write_7_stage_43;
      dark_dark_update_0_write_write_7_stage_45 <= dark_dark_update_0_write_write_7_stage_44;
      dark_dark_update_0_write_write_7_stage_46 <= dark_dark_update_0_write_write_7_stage_45;
      dark_dark_update_0_write_write_7_stage_47 <= dark_dark_update_0_write_write_7_stage_46;
      dark_dark_update_0_write_write_7_stage_48 <= dark_dark_update_0_write_write_7_stage_47;
      dark_dark_update_0_write_write_7_stage_49 <= dark_dark_update_0_write_write_7_stage_48;
      dark_dark_update_0_write_write_7_stage_50 <= dark_dark_update_0_write_write_7_stage_49;
      dark_dark_update_0_write_write_7_stage_51 <= dark_dark_update_0_write_write_7_stage_50;
      dark_dark_update_0_write_write_7_stage_52 <= dark_dark_update_0_write_write_7_stage_51;
      dark_dark_update_0_write_write_7_stage_53 <= dark_dark_update_0_write_write_7_stage_52;
      dark_dark_update_0_write_write_7_stage_54 <= dark_dark_update_0_write_write_7_stage_53;
      dark_dark_update_0_write_write_7_stage_55 <= dark_dark_update_0_write_write_7_stage_54;
      dark_dark_update_0_write_write_7_stage_56 <= dark_dark_update_0_write_write_7_stage_55;
      dark_dark_update_0_write_write_7_stage_57 <= dark_dark_update_0_write_write_7_stage_56;
      dark_dark_update_0_write_write_7_stage_58 <= dark_dark_update_0_write_write_7_stage_57;
      dark_dark_update_0_write_write_7_stage_59 <= dark_dark_update_0_write_write_7_stage_58;
      dark_dark_update_0_write_write_7_stage_60 <= dark_dark_update_0_write_write_7_stage_59;
      dark_dark_update_0_write_write_7_stage_61 <= dark_dark_update_0_write_write_7_stage_60;
      dark_dark_update_0_write_write_7_stage_62 <= dark_dark_update_0_write_write_7_stage_61;
      dark_dark_update_0_write_write_7_stage_63 <= dark_dark_update_0_write_write_7_stage_62;
      dark_dark_update_0_write_write_7_stage_64 <= dark_dark_update_0_write_write_7_stage_63;
      dark_dark_update_0_write_write_7_stage_65 <= dark_dark_update_0_write_write_7_stage_64;
      dark_dark_update_0_write_write_7_stage_66 <= dark_dark_update_0_write_write_7_stage_65;
      dark_dark_update_0_write_write_7_stage_67 <= dark_dark_update_0_write_write_7_stage_66;
      dark_dark_update_0_write_write_7_stage_68 <= dark_dark_update_0_write_write_7_stage_67;
      dark_dark_update_0_write_write_7_stage_69 <= dark_dark_update_0_write_write_7_stage_68;
      dark_dark_update_0_write_write_7_stage_70 <= dark_dark_update_0_write_write_7_stage_69;
      dark_dark_update_0_write_write_7_stage_71 <= dark_dark_update_0_write_write_7_stage_70;
      dark_dark_update_0_write_write_7_stage_72 <= dark_dark_update_0_write_write_7_stage_71;
      dark_dark_update_0_write_write_7_stage_73 <= dark_dark_update_0_write_write_7_stage_72;
      dark_dark_update_0_write_write_7_stage_74 <= dark_dark_update_0_write_write_7_stage_73;
      dark_dark_update_0_write_write_7_stage_75 <= dark_dark_update_0_write_write_7_stage_74;
      dark_dark_update_0_write_write_7_stage_76 <= dark_dark_update_0_write_write_7_stage_75;
      dark_dark_update_0_write_write_7_stage_77 <= dark_dark_update_0_write_write_7_stage_76;
      dark_dark_update_0_write_write_7_stage_78 <= dark_dark_update_0_write_write_7_stage_77;
      dark_dark_update_0_write_write_7_stage_79 <= dark_dark_update_0_write_write_7_stage_78;
      dark_dark_update_0_write_write_7_stage_80 <= dark_dark_update_0_write_write_7_stage_79;
      dark_dark_update_0_write_write_7_stage_81 <= dark_dark_update_0_write_write_7_stage_80;
      dark_dark_update_0_write_write_7_stage_82 <= dark_dark_update_0_write_write_7_stage_81;
      dark_dark_update_0_write_write_7_stage_83 <= dark_dark_update_0_write_write_7_stage_82;
      dark_dark_update_0_write_write_7_stage_84 <= dark_dark_update_0_write_write_7_stage_83;
      dark_dark_update_0_write_write_7_stage_85 <= dark_dark_update_0_write_write_7_stage_84;
      dark_dark_update_0_write_write_7_stage_86 <= dark_dark_update_0_write_write_7_stage_85;
      dark_dark_update_0_write_write_7_stage_87 <= dark_dark_update_0_write_write_7_stage_86;
      dark_dark_update_0_write_write_7_stage_88 <= dark_dark_update_0_write_write_7_stage_87;
      dark_dark_update_0_write_write_7_stage_89 <= dark_dark_update_0_write_write_7_stage_88;
      dark_dark_update_0_write_write_7_stage_90 <= dark_dark_update_0_write_write_7_stage_89;
      dark_dark_update_0_write_write_7_stage_91 <= dark_dark_update_0_write_write_7_stage_90;
      dark_dark_update_0_write_write_7_stage_92 <= dark_dark_update_0_write_write_7_stage_91;
      dark_dark_update_0_write_write_7_stage_93 <= dark_dark_update_0_write_write_7_stage_92;
      dark_dark_update_0_write_write_7_stage_94 <= dark_dark_update_0_write_write_7_stage_93;
      dark_dark_update_0_write_write_7_stage_95 <= dark_dark_update_0_write_write_7_stage_94;
      dark_dark_update_0_write_write_7_stage_96 <= dark_dark_update_0_write_write_7_stage_95;
      dark_dark_update_0_write_write_7_stage_97 <= dark_dark_update_0_write_write_7_stage_96;
      dark_dark_update_0_write_write_7_stage_98 <= dark_dark_update_0_write_write_7_stage_97;
      dark_dark_update_0_write_write_7_stage_99 <= dark_dark_update_0_write_write_7_stage_98;
      dark_dark_update_0_write_write_7_stage_100 <= dark_dark_update_0_write_write_7_stage_99;
      dark_dark_update_0_write_write_7_stage_101 <= dark_dark_update_0_write_write_7_stage_100;
      dark_dark_update_0_write_write_7_stage_102 <= dark_dark_update_0_write_write_7_stage_101;
      dark_dark_update_0_write_write_7_stage_103 <= dark_dark_update_0_write_write_7_stage_102;
      dark_dark_update_0_write_write_7_stage_104 <= dark_dark_update_0_write_write_7_stage_103;
      dark_dark_update_0_write_write_7_stage_105 <= dark_dark_update_0_write_write_7_stage_104;
      dark_dark_update_0_write_write_7_stage_106 <= dark_dark_update_0_write_write_7_stage_105;
      dark_dark_update_0_write_write_7_stage_107 <= dark_dark_update_0_write_write_7_stage_106;
      dark_dark_update_0_write_write_7_stage_108 <= dark_dark_update_0_write_write_7_stage_107;
      dark_dark_update_0_write_write_7_stage_109 <= dark_dark_update_0_write_write_7_stage_108;
      dark_dark_update_0_write_write_7_stage_110 <= dark_dark_update_0_write_write_7_stage_109;
      dark_dark_update_0_write_write_7_stage_111 <= dark_dark_update_0_write_write_7_stage_110;
      dark_dark_update_0_write_write_7_stage_112 <= dark_dark_update_0_write_write_7_stage_111;
      dark_dark_update_0_write_write_7_stage_113 <= dark_dark_update_0_write_write_7_stage_112;
      dark_dark_update_0_write_write_7_stage_114 <= dark_dark_update_0_write_write_7_stage_113;
      dark_dark_update_0_write_write_7_stage_115 <= dark_dark_update_0_write_write_7_stage_114;
      dark_dark_update_0_write_write_7_stage_116 <= dark_dark_update_0_write_write_7_stage_115;
      dark_dark_update_0_write_write_7_stage_117 <= dark_dark_update_0_write_write_7_stage_116;
      dark_dark_update_0_write_write_7_stage_118 <= dark_dark_update_0_write_write_7_stage_117;
      dark_dark_update_0_write_write_7_stage_119 <= dark_dark_update_0_write_write_7_stage_118;
      dark_dark_update_0_write_write_7_stage_120 <= dark_dark_update_0_write_write_7_stage_119;
      dark_dark_update_0_write_write_7_stage_121 <= dark_dark_update_0_write_write_7_stage_120;
      dark_dark_update_0_write_write_7_stage_122 <= dark_dark_update_0_write_write_7_stage_121;
      dark_dark_update_0_write_write_7_stage_123 <= dark_dark_update_0_write_write_7_stage_122;
      dark_dark_update_0_write_write_7_stage_124 <= dark_dark_update_0_write_write_7_stage_123;
      dark_dark_update_0_write_write_7_stage_125 <= dark_dark_update_0_write_write_7_stage_124;
      dark_dark_update_0_write_write_7_stage_126 <= dark_dark_update_0_write_write_7_stage_125;
      dark_dark_update_0_write_write_7_stage_127 <= dark_dark_update_0_write_write_7_stage_126;
      dark_dark_update_0_write_write_7_stage_128 <= dark_dark_update_0_write_write_7_stage_127;
      dark_dark_update_0_write_write_7_stage_129 <= dark_dark_update_0_write_write_7_stage_128;
      dark_dark_update_0_write_write_7_stage_130 <= dark_dark_update_0_write_write_7_stage_129;
      dark_dark_update_0_write_write_7_stage_131 <= dark_dark_update_0_write_write_7_stage_130;
      dark_dark_update_0_write_write_7_stage_132 <= dark_dark_update_0_write_write_7_stage_131;
      dark_dark_update_0_write_write_7_stage_133 <= dark_dark_update_0_write_write_7_stage_132;
      dark_dark_update_0_write_write_7_stage_134 <= dark_dark_update_0_write_write_7_stage_133;
      dark_dark_update_0_write_write_7_stage_135 <= dark_dark_update_0_write_write_7_stage_134;
      dark_dark_update_0_write_write_7_stage_136 <= dark_dark_update_0_write_write_7_stage_135;
      dark_dark_update_0_write_write_7_stage_137 <= dark_dark_update_0_write_write_7_stage_136;
      dark_dark_update_0_write_write_7_stage_138 <= dark_dark_update_0_write_write_7_stage_137;
      dark_dark_update_0_write_write_7_stage_139 <= dark_dark_update_0_write_write_7_stage_138;
      dark_dark_update_0_write_write_7_stage_140 <= dark_dark_update_0_write_write_7_stage_139;
      dark_dark_update_0_write_write_7_stage_141 <= dark_dark_update_0_write_write_7_stage_140;
      dark_dark_update_0_write_write_7_stage_142 <= dark_dark_update_0_write_write_7_stage_141;
      dark_dark_update_0_write_write_7_stage_143 <= dark_dark_update_0_write_write_7_stage_142;
      dark_dark_update_0_write_write_7_stage_144 <= dark_dark_update_0_write_write_7_stage_143;
      dark_dark_update_0_write_write_7_stage_145 <= dark_dark_update_0_write_write_7_stage_144;
      dark_dark_update_0_write_write_7_stage_146 <= dark_dark_update_0_write_write_7_stage_145;
      dark_dark_update_0_write_write_7_stage_147 <= dark_dark_update_0_write_write_7_stage_146;
      dark_dark_update_0_write_write_7_stage_148 <= dark_dark_update_0_write_write_7_stage_147;
      dark_dark_update_0_write_write_7_stage_149 <= dark_dark_update_0_write_write_7_stage_148;
      dark_dark_update_0_write_write_7_stage_150 <= dark_dark_update_0_write_write_7_stage_149;
      dark_dark_update_0_write_write_7_stage_151 <= dark_dark_update_0_write_write_7_stage_150;
      dark_dark_update_0_write_write_7_stage_152 <= dark_dark_update_0_write_write_7_stage_151;
      dark_dark_update_0_write_write_7_stage_153 <= dark_dark_update_0_write_write_7_stage_152;
      dark_dark_update_0_write_write_7_stage_154 <= dark_dark_update_0_write_write_7_stage_153;
      dark_dark_update_0_write_write_7_stage_155 <= dark_dark_update_0_write_write_7_stage_154;
      dark_dark_update_0_write_write_7_stage_156 <= dark_dark_update_0_write_write_7_stage_155;
      dark_dark_update_0_write_write_7_stage_157 <= dark_dark_update_0_write_write_7_stage_156;
      dark_dark_update_0_write_write_7_stage_158 <= dark_dark_update_0_write_write_7_stage_157;
      dark_dark_update_0_write_write_7_stage_159 <= dark_dark_update_0_write_write_7_stage_158;
      dark_dark_update_0_write_write_7_stage_160 <= dark_dark_update_0_write_write_7_stage_159;
      dark_dark_update_0_write_write_7_stage_161 <= dark_dark_update_0_write_write_7_stage_160;
      dark_dark_update_0_write_write_7_stage_162 <= dark_dark_update_0_write_write_7_stage_161;
      dark_dark_update_0_write_write_7_stage_163 <= dark_dark_update_0_write_write_7_stage_162;
      dark_dark_update_0_write_write_7_stage_164 <= dark_dark_update_0_write_write_7_stage_163;
      dark_dark_update_0_write_write_7_stage_165 <= dark_dark_update_0_write_write_7_stage_164;
      dark_dark_update_0_write_write_7_stage_166 <= dark_dark_update_0_write_write_7_stage_165;
      dark_dark_update_0_write_write_7_stage_167 <= dark_dark_update_0_write_write_7_stage_166;
      dark_dark_update_0_write_write_7_stage_168 <= dark_dark_update_0_write_write_7_stage_167;
      dark_dark_update_0_write_write_7_stage_169 <= dark_dark_update_0_write_write_7_stage_168;
      dark_dark_update_0_write_write_7_stage_170 <= dark_dark_update_0_write_write_7_stage_169;
      dark_dark_update_0_write_write_7_stage_171 <= dark_dark_update_0_write_write_7_stage_170;
      dark_dark_update_0_write_write_7_stage_172 <= dark_dark_update_0_write_write_7_stage_171;
      dark_dark_update_0_write_write_7_stage_173 <= dark_dark_update_0_write_write_7_stage_172;
      dark_dark_update_0_write_write_7_stage_174 <= dark_dark_update_0_write_write_7_stage_173;
      dark_dark_update_0_write_write_7_stage_175 <= dark_dark_update_0_write_write_7_stage_174;
      dark_dark_update_0_write_write_7_stage_176 <= dark_dark_update_0_write_write_7_stage_175;
      dark_dark_update_0_write_write_7_stage_177 <= dark_dark_update_0_write_write_7_stage_176;
      dark_dark_update_0_write_write_7_stage_178 <= dark_dark_update_0_write_write_7_stage_177;
      dark_dark_update_0_write_write_7_stage_179 <= dark_dark_update_0_write_write_7_stage_178;
      dark_dark_update_0_write_write_7_stage_180 <= dark_dark_update_0_write_write_7_stage_179;
      dark_dark_update_0_write_write_7_stage_181 <= dark_dark_update_0_write_write_7_stage_180;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_17 <= dark_dark_gauss_blur_1_update_0_read_read_10;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_18 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_17;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_19 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_18;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_20 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_19;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_21 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_20;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_22 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_21;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_23 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_22;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_24 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_23;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_25 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_24;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_26 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_25;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_27 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_26;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_28 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_27;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_29 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_28;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_30 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_29;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_31 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_30;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_32 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_31;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_33 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_32;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_34 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_33;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_35 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_34;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_36 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_35;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_37 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_36;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_38 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_37;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_39 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_38;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_40 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_39;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_41 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_40;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_42 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_41;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_43 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_42;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_44 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_43;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_45 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_44;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_46 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_45;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_47 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_46;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_48 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_47;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_49 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_48;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_50 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_49;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_51 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_50;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_52 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_51;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_53 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_52;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_54 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_53;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_55 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_54;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_56 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_55;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_57 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_56;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_58 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_57;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_59 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_58;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_60 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_59;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_61 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_60;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_62 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_61;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_63 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_62;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_64 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_63;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_65 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_64;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_66 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_65;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_67 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_66;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_68 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_67;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_69 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_68;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_70 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_69;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_71 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_70;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_72 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_71;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_73 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_72;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_74 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_73;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_75 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_74;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_76 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_75;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_77 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_76;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_78 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_77;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_79 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_78;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_80 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_79;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_81 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_80;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_82 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_81;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_83 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_82;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_84 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_83;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_85 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_84;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_86 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_85;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_87 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_86;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_88 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_87;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_89 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_88;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_90 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_89;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_91 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_90;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_92 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_91;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_93 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_92;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_94 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_93;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_95 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_94;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_96 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_95;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_97 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_96;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_98 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_97;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_99 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_98;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_100 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_99;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_101 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_100;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_102 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_101;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_103 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_102;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_104 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_103;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_105 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_104;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_106 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_105;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_107 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_106;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_108 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_107;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_109 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_108;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_110 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_109;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_111 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_110;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_112 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_111;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_113 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_112;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_114 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_113;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_115 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_114;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_116 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_115;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_117 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_116;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_118 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_117;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_119 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_118;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_120 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_119;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_121 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_120;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_122 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_121;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_123 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_122;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_124 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_123;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_125 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_124;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_126 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_125;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_127 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_126;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_128 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_127;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_129 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_128;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_130 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_129;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_131 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_130;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_132 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_131;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_133 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_132;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_134 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_133;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_135 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_134;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_136 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_135;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_137 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_136;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_138 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_137;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_139 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_138;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_140 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_139;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_141 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_140;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_142 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_141;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_143 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_142;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_144 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_143;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_145 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_144;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_146 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_145;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_147 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_146;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_148 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_147;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_149 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_148;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_150 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_149;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_151 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_150;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_152 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_151;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_153 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_152;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_154 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_153;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_155 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_154;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_156 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_155;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_157 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_156;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_158 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_157;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_159 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_158;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_160 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_159;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_161 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_160;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_162 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_161;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_163 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_162;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_164 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_163;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_165 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_164;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_166 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_165;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_167 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_166;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_168 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_167;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_169 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_168;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_170 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_169;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_171 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_170;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_172 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_171;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_173 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_172;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_174 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_173;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_175 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_174;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_176 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_175;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_177 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_176;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_178 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_177;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_179 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_178;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_180 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_179;
      dark_dark_gauss_blur_1_update_0_read_read_10_stage_181 <= dark_dark_gauss_blur_1_update_0_read_read_10_stage_180;
      dark_gauss_blur_1_update_0_stage_18 <= dark_gauss_blur_1_update_0;
      dark_gauss_blur_1_update_0_stage_19 <= dark_gauss_blur_1_update_0_stage_18;
      dark_gauss_blur_1_update_0_stage_20 <= dark_gauss_blur_1_update_0_stage_19;
      dark_gauss_blur_1_update_0_stage_21 <= dark_gauss_blur_1_update_0_stage_20;
      dark_gauss_blur_1_update_0_stage_22 <= dark_gauss_blur_1_update_0_stage_21;
      dark_gauss_blur_1_update_0_stage_23 <= dark_gauss_blur_1_update_0_stage_22;
      dark_gauss_blur_1_update_0_stage_24 <= dark_gauss_blur_1_update_0_stage_23;
      dark_gauss_blur_1_update_0_stage_25 <= dark_gauss_blur_1_update_0_stage_24;
      dark_gauss_blur_1_update_0_stage_26 <= dark_gauss_blur_1_update_0_stage_25;
      dark_gauss_blur_1_update_0_stage_27 <= dark_gauss_blur_1_update_0_stage_26;
      dark_gauss_blur_1_update_0_stage_28 <= dark_gauss_blur_1_update_0_stage_27;
      dark_gauss_blur_1_update_0_stage_29 <= dark_gauss_blur_1_update_0_stage_28;
      dark_gauss_blur_1_update_0_stage_30 <= dark_gauss_blur_1_update_0_stage_29;
      dark_gauss_blur_1_update_0_stage_31 <= dark_gauss_blur_1_update_0_stage_30;
      dark_gauss_blur_1_update_0_stage_32 <= dark_gauss_blur_1_update_0_stage_31;
      dark_gauss_blur_1_update_0_stage_33 <= dark_gauss_blur_1_update_0_stage_32;
      dark_gauss_blur_1_update_0_stage_34 <= dark_gauss_blur_1_update_0_stage_33;
      dark_gauss_blur_1_update_0_stage_35 <= dark_gauss_blur_1_update_0_stage_34;
      dark_gauss_blur_1_update_0_stage_36 <= dark_gauss_blur_1_update_0_stage_35;
      dark_gauss_blur_1_update_0_stage_37 <= dark_gauss_blur_1_update_0_stage_36;
      dark_gauss_blur_1_update_0_stage_38 <= dark_gauss_blur_1_update_0_stage_37;
      dark_gauss_blur_1_update_0_stage_39 <= dark_gauss_blur_1_update_0_stage_38;
      dark_gauss_blur_1_update_0_stage_40 <= dark_gauss_blur_1_update_0_stage_39;
      dark_gauss_blur_1_update_0_stage_41 <= dark_gauss_blur_1_update_0_stage_40;
      dark_gauss_blur_1_update_0_stage_42 <= dark_gauss_blur_1_update_0_stage_41;
      dark_gauss_blur_1_update_0_stage_43 <= dark_gauss_blur_1_update_0_stage_42;
      dark_gauss_blur_1_update_0_stage_44 <= dark_gauss_blur_1_update_0_stage_43;
      dark_gauss_blur_1_update_0_stage_45 <= dark_gauss_blur_1_update_0_stage_44;
      dark_gauss_blur_1_update_0_stage_46 <= dark_gauss_blur_1_update_0_stage_45;
      dark_gauss_blur_1_update_0_stage_47 <= dark_gauss_blur_1_update_0_stage_46;
      dark_gauss_blur_1_update_0_stage_48 <= dark_gauss_blur_1_update_0_stage_47;
      dark_gauss_blur_1_update_0_stage_49 <= dark_gauss_blur_1_update_0_stage_48;
      dark_gauss_blur_1_update_0_stage_50 <= dark_gauss_blur_1_update_0_stage_49;
      dark_gauss_blur_1_update_0_stage_51 <= dark_gauss_blur_1_update_0_stage_50;
      dark_gauss_blur_1_update_0_stage_52 <= dark_gauss_blur_1_update_0_stage_51;
      dark_gauss_blur_1_update_0_stage_53 <= dark_gauss_blur_1_update_0_stage_52;
      dark_gauss_blur_1_update_0_stage_54 <= dark_gauss_blur_1_update_0_stage_53;
      dark_gauss_blur_1_update_0_stage_55 <= dark_gauss_blur_1_update_0_stage_54;
      dark_gauss_blur_1_update_0_stage_56 <= dark_gauss_blur_1_update_0_stage_55;
      dark_gauss_blur_1_update_0_stage_57 <= dark_gauss_blur_1_update_0_stage_56;
      dark_gauss_blur_1_update_0_stage_58 <= dark_gauss_blur_1_update_0_stage_57;
      dark_gauss_blur_1_update_0_stage_59 <= dark_gauss_blur_1_update_0_stage_58;
      dark_gauss_blur_1_update_0_stage_60 <= dark_gauss_blur_1_update_0_stage_59;
      dark_gauss_blur_1_update_0_stage_61 <= dark_gauss_blur_1_update_0_stage_60;
      dark_gauss_blur_1_update_0_stage_62 <= dark_gauss_blur_1_update_0_stage_61;
      dark_gauss_blur_1_update_0_stage_63 <= dark_gauss_blur_1_update_0_stage_62;
      dark_gauss_blur_1_update_0_stage_64 <= dark_gauss_blur_1_update_0_stage_63;
      dark_gauss_blur_1_update_0_stage_65 <= dark_gauss_blur_1_update_0_stage_64;
      dark_gauss_blur_1_update_0_stage_66 <= dark_gauss_blur_1_update_0_stage_65;
      dark_gauss_blur_1_update_0_stage_67 <= dark_gauss_blur_1_update_0_stage_66;
      dark_gauss_blur_1_update_0_stage_68 <= dark_gauss_blur_1_update_0_stage_67;
      dark_gauss_blur_1_update_0_stage_69 <= dark_gauss_blur_1_update_0_stage_68;
      dark_gauss_blur_1_update_0_stage_70 <= dark_gauss_blur_1_update_0_stage_69;
      dark_gauss_blur_1_update_0_stage_71 <= dark_gauss_blur_1_update_0_stage_70;
      dark_gauss_blur_1_update_0_stage_72 <= dark_gauss_blur_1_update_0_stage_71;
      dark_gauss_blur_1_update_0_stage_73 <= dark_gauss_blur_1_update_0_stage_72;
      dark_gauss_blur_1_update_0_stage_74 <= dark_gauss_blur_1_update_0_stage_73;
      dark_gauss_blur_1_update_0_stage_75 <= dark_gauss_blur_1_update_0_stage_74;
      dark_gauss_blur_1_update_0_stage_76 <= dark_gauss_blur_1_update_0_stage_75;
      dark_gauss_blur_1_update_0_stage_77 <= dark_gauss_blur_1_update_0_stage_76;
      dark_gauss_blur_1_update_0_stage_78 <= dark_gauss_blur_1_update_0_stage_77;
      dark_gauss_blur_1_update_0_stage_79 <= dark_gauss_blur_1_update_0_stage_78;
      dark_gauss_blur_1_update_0_stage_80 <= dark_gauss_blur_1_update_0_stage_79;
      dark_gauss_blur_1_update_0_stage_81 <= dark_gauss_blur_1_update_0_stage_80;
      dark_gauss_blur_1_update_0_stage_82 <= dark_gauss_blur_1_update_0_stage_81;
      dark_gauss_blur_1_update_0_stage_83 <= dark_gauss_blur_1_update_0_stage_82;
      dark_gauss_blur_1_update_0_stage_84 <= dark_gauss_blur_1_update_0_stage_83;
      dark_gauss_blur_1_update_0_stage_85 <= dark_gauss_blur_1_update_0_stage_84;
      dark_gauss_blur_1_update_0_stage_86 <= dark_gauss_blur_1_update_0_stage_85;
      dark_gauss_blur_1_update_0_stage_87 <= dark_gauss_blur_1_update_0_stage_86;
      dark_gauss_blur_1_update_0_stage_88 <= dark_gauss_blur_1_update_0_stage_87;
      dark_gauss_blur_1_update_0_stage_89 <= dark_gauss_blur_1_update_0_stage_88;
      dark_gauss_blur_1_update_0_stage_90 <= dark_gauss_blur_1_update_0_stage_89;
      dark_gauss_blur_1_update_0_stage_91 <= dark_gauss_blur_1_update_0_stage_90;
      dark_gauss_blur_1_update_0_stage_92 <= dark_gauss_blur_1_update_0_stage_91;
      dark_gauss_blur_1_update_0_stage_93 <= dark_gauss_blur_1_update_0_stage_92;
      dark_gauss_blur_1_update_0_stage_94 <= dark_gauss_blur_1_update_0_stage_93;
      dark_gauss_blur_1_update_0_stage_95 <= dark_gauss_blur_1_update_0_stage_94;
      dark_gauss_blur_1_update_0_stage_96 <= dark_gauss_blur_1_update_0_stage_95;
      dark_gauss_blur_1_update_0_stage_97 <= dark_gauss_blur_1_update_0_stage_96;
      dark_gauss_blur_1_update_0_stage_98 <= dark_gauss_blur_1_update_0_stage_97;
      dark_gauss_blur_1_update_0_stage_99 <= dark_gauss_blur_1_update_0_stage_98;
      dark_gauss_blur_1_update_0_stage_100 <= dark_gauss_blur_1_update_0_stage_99;
      dark_gauss_blur_1_update_0_stage_101 <= dark_gauss_blur_1_update_0_stage_100;
      dark_gauss_blur_1_update_0_stage_102 <= dark_gauss_blur_1_update_0_stage_101;
      dark_gauss_blur_1_update_0_stage_103 <= dark_gauss_blur_1_update_0_stage_102;
      dark_gauss_blur_1_update_0_stage_104 <= dark_gauss_blur_1_update_0_stage_103;
      dark_gauss_blur_1_update_0_stage_105 <= dark_gauss_blur_1_update_0_stage_104;
      dark_gauss_blur_1_update_0_stage_106 <= dark_gauss_blur_1_update_0_stage_105;
      dark_gauss_blur_1_update_0_stage_107 <= dark_gauss_blur_1_update_0_stage_106;
      dark_gauss_blur_1_update_0_stage_108 <= dark_gauss_blur_1_update_0_stage_107;
      dark_gauss_blur_1_update_0_stage_109 <= dark_gauss_blur_1_update_0_stage_108;
      dark_gauss_blur_1_update_0_stage_110 <= dark_gauss_blur_1_update_0_stage_109;
      dark_gauss_blur_1_update_0_stage_111 <= dark_gauss_blur_1_update_0_stage_110;
      dark_gauss_blur_1_update_0_stage_112 <= dark_gauss_blur_1_update_0_stage_111;
      dark_gauss_blur_1_update_0_stage_113 <= dark_gauss_blur_1_update_0_stage_112;
      dark_gauss_blur_1_update_0_stage_114 <= dark_gauss_blur_1_update_0_stage_113;
      dark_gauss_blur_1_update_0_stage_115 <= dark_gauss_blur_1_update_0_stage_114;
      dark_gauss_blur_1_update_0_stage_116 <= dark_gauss_blur_1_update_0_stage_115;
      dark_gauss_blur_1_update_0_stage_117 <= dark_gauss_blur_1_update_0_stage_116;
      dark_gauss_blur_1_update_0_stage_118 <= dark_gauss_blur_1_update_0_stage_117;
      dark_gauss_blur_1_update_0_stage_119 <= dark_gauss_blur_1_update_0_stage_118;
      dark_gauss_blur_1_update_0_stage_120 <= dark_gauss_blur_1_update_0_stage_119;
      dark_gauss_blur_1_update_0_stage_121 <= dark_gauss_blur_1_update_0_stage_120;
      dark_gauss_blur_1_update_0_stage_122 <= dark_gauss_blur_1_update_0_stage_121;
      dark_gauss_blur_1_update_0_stage_123 <= dark_gauss_blur_1_update_0_stage_122;
      dark_gauss_blur_1_update_0_stage_124 <= dark_gauss_blur_1_update_0_stage_123;
      dark_gauss_blur_1_update_0_stage_125 <= dark_gauss_blur_1_update_0_stage_124;
      dark_gauss_blur_1_update_0_stage_126 <= dark_gauss_blur_1_update_0_stage_125;
      dark_gauss_blur_1_update_0_stage_127 <= dark_gauss_blur_1_update_0_stage_126;
      dark_gauss_blur_1_update_0_stage_128 <= dark_gauss_blur_1_update_0_stage_127;
      dark_gauss_blur_1_update_0_stage_129 <= dark_gauss_blur_1_update_0_stage_128;
      dark_gauss_blur_1_update_0_stage_130 <= dark_gauss_blur_1_update_0_stage_129;
      dark_gauss_blur_1_update_0_stage_131 <= dark_gauss_blur_1_update_0_stage_130;
      dark_gauss_blur_1_update_0_stage_132 <= dark_gauss_blur_1_update_0_stage_131;
      dark_gauss_blur_1_update_0_stage_133 <= dark_gauss_blur_1_update_0_stage_132;
      dark_gauss_blur_1_update_0_stage_134 <= dark_gauss_blur_1_update_0_stage_133;
      dark_gauss_blur_1_update_0_stage_135 <= dark_gauss_blur_1_update_0_stage_134;
      dark_gauss_blur_1_update_0_stage_136 <= dark_gauss_blur_1_update_0_stage_135;
      dark_gauss_blur_1_update_0_stage_137 <= dark_gauss_blur_1_update_0_stage_136;
      dark_gauss_blur_1_update_0_stage_138 <= dark_gauss_blur_1_update_0_stage_137;
      dark_gauss_blur_1_update_0_stage_139 <= dark_gauss_blur_1_update_0_stage_138;
      dark_gauss_blur_1_update_0_stage_140 <= dark_gauss_blur_1_update_0_stage_139;
      dark_gauss_blur_1_update_0_stage_141 <= dark_gauss_blur_1_update_0_stage_140;
      dark_gauss_blur_1_update_0_stage_142 <= dark_gauss_blur_1_update_0_stage_141;
      dark_gauss_blur_1_update_0_stage_143 <= dark_gauss_blur_1_update_0_stage_142;
      dark_gauss_blur_1_update_0_stage_144 <= dark_gauss_blur_1_update_0_stage_143;
      dark_gauss_blur_1_update_0_stage_145 <= dark_gauss_blur_1_update_0_stage_144;
      dark_gauss_blur_1_update_0_stage_146 <= dark_gauss_blur_1_update_0_stage_145;
      dark_gauss_blur_1_update_0_stage_147 <= dark_gauss_blur_1_update_0_stage_146;
      dark_gauss_blur_1_update_0_stage_148 <= dark_gauss_blur_1_update_0_stage_147;
      dark_gauss_blur_1_update_0_stage_149 <= dark_gauss_blur_1_update_0_stage_148;
      dark_gauss_blur_1_update_0_stage_150 <= dark_gauss_blur_1_update_0_stage_149;
      dark_gauss_blur_1_update_0_stage_151 <= dark_gauss_blur_1_update_0_stage_150;
      dark_gauss_blur_1_update_0_stage_152 <= dark_gauss_blur_1_update_0_stage_151;
      dark_gauss_blur_1_update_0_stage_153 <= dark_gauss_blur_1_update_0_stage_152;
      dark_gauss_blur_1_update_0_stage_154 <= dark_gauss_blur_1_update_0_stage_153;
      dark_gauss_blur_1_update_0_stage_155 <= dark_gauss_blur_1_update_0_stage_154;
      dark_gauss_blur_1_update_0_stage_156 <= dark_gauss_blur_1_update_0_stage_155;
      dark_gauss_blur_1_update_0_stage_157 <= dark_gauss_blur_1_update_0_stage_156;
      dark_gauss_blur_1_update_0_stage_158 <= dark_gauss_blur_1_update_0_stage_157;
      dark_gauss_blur_1_update_0_stage_159 <= dark_gauss_blur_1_update_0_stage_158;
      dark_gauss_blur_1_update_0_stage_160 <= dark_gauss_blur_1_update_0_stage_159;
      dark_gauss_blur_1_update_0_stage_161 <= dark_gauss_blur_1_update_0_stage_160;
      dark_gauss_blur_1_update_0_stage_162 <= dark_gauss_blur_1_update_0_stage_161;
      dark_gauss_blur_1_update_0_stage_163 <= dark_gauss_blur_1_update_0_stage_162;
      dark_gauss_blur_1_update_0_stage_164 <= dark_gauss_blur_1_update_0_stage_163;
      dark_gauss_blur_1_update_0_stage_165 <= dark_gauss_blur_1_update_0_stage_164;
      dark_gauss_blur_1_update_0_stage_166 <= dark_gauss_blur_1_update_0_stage_165;
      dark_gauss_blur_1_update_0_stage_167 <= dark_gauss_blur_1_update_0_stage_166;
      dark_gauss_blur_1_update_0_stage_168 <= dark_gauss_blur_1_update_0_stage_167;
      dark_gauss_blur_1_update_0_stage_169 <= dark_gauss_blur_1_update_0_stage_168;
      dark_gauss_blur_1_update_0_stage_170 <= dark_gauss_blur_1_update_0_stage_169;
      dark_gauss_blur_1_update_0_stage_171 <= dark_gauss_blur_1_update_0_stage_170;
      dark_gauss_blur_1_update_0_stage_172 <= dark_gauss_blur_1_update_0_stage_171;
      dark_gauss_blur_1_update_0_stage_173 <= dark_gauss_blur_1_update_0_stage_172;
      dark_gauss_blur_1_update_0_stage_174 <= dark_gauss_blur_1_update_0_stage_173;
      dark_gauss_blur_1_update_0_stage_175 <= dark_gauss_blur_1_update_0_stage_174;
      dark_gauss_blur_1_update_0_stage_176 <= dark_gauss_blur_1_update_0_stage_175;
      dark_gauss_blur_1_update_0_stage_177 <= dark_gauss_blur_1_update_0_stage_176;
      dark_gauss_blur_1_update_0_stage_178 <= dark_gauss_blur_1_update_0_stage_177;
      dark_gauss_blur_1_update_0_stage_179 <= dark_gauss_blur_1_update_0_stage_178;
      dark_gauss_blur_1_update_0_stage_180 <= dark_gauss_blur_1_update_0_stage_179;
      dark_gauss_blur_1_update_0_stage_181 <= dark_gauss_blur_1_update_0_stage_180;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_60 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_61 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_60;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_62 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_61;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_63 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_62;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_64 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_63;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_65 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_64;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_66 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_65;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_67 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_66;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_68 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_67;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_69 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_68;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_70 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_69;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_71 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_70;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_72 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_71;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_73 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_72;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_74 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_73;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_75 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_74;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_76 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_75;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_77 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_76;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_78 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_77;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_79 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_78;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_80 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_79;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_81 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_80;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_82 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_81;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_83 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_82;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_84 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_83;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_85 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_84;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_86 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_85;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_87 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_86;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_88 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_87;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_89 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_88;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_90 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_89;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_91 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_90;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_92 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_91;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_93 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_92;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_94 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_93;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_95 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_94;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_96 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_95;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_97 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_96;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_98 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_97;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_99 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_98;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_100 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_99;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_101 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_100;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_102 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_101;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_103 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_102;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_104 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_103;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_105 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_104;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_106 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_105;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_107 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_106;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_108 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_107;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_109 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_108;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_110 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_109;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_111 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_110;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_112 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_111;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_113 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_112;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_114 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_113;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_115 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_114;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_116 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_115;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_117 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_116;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_118 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_117;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_119 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_118;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_120 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_119;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_121 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_120;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_122 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_121;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_123 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_122;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_124 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_123;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_125 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_124;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_126 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_125;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_127 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_126;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_128 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_127;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_129 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_128;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_130 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_129;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_131 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_130;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_132 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_131;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_133 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_132;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_134 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_133;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_135 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_134;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_136 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_135;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_137 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_136;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_138 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_137;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_139 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_138;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_140 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_139;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_141 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_140;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_142 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_141;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_143 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_142;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_144 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_143;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_145 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_144;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_146 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_145;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_147 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_146;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_148 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_147;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_149 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_148;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_150 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_149;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_151 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_150;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_152 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_151;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_153 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_152;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_154 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_153;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_155 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_154;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_156 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_155;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_157 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_156;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_158 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_157;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_159 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_158;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_160 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_159;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_161 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_160;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_162 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_161;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_163 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_162;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_164 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_163;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_165 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_164;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_166 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_165;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_167 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_166;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_168 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_167;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_169 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_168;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_170 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_169;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_171 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_170;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_172 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_171;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_173 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_172;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_174 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_173;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_175 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_174;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_176 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_175;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_177 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_176;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_178 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_177;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_179 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_178;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_180 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_179;
      bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_181 <= bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39_stage_180;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_19 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_20 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_19;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_21 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_20;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_22 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_21;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_23 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_22;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_24 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_23;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_25 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_24;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_26 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_25;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_27 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_26;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_28 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_27;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_29 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_28;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_30 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_29;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_31 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_30;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_32 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_31;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_33 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_32;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_34 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_33;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_35 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_34;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_36 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_35;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_37 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_36;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_38 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_37;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_39 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_38;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_40 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_39;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_41 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_40;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_42 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_41;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_43 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_42;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_44 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_43;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_45 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_44;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_46 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_45;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_47 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_46;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_48 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_47;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_49 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_48;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_50 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_49;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_51 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_50;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_52 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_51;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_53 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_52;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_54 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_53;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_55 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_54;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_56 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_55;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_57 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_56;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_58 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_57;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_59 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_58;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_60 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_59;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_61 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_60;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_62 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_61;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_63 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_62;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_64 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_63;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_65 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_64;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_66 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_65;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_67 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_66;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_68 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_67;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_69 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_68;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_70 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_69;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_71 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_70;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_72 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_71;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_73 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_72;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_74 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_73;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_75 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_74;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_76 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_75;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_77 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_76;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_78 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_77;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_79 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_78;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_80 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_79;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_81 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_80;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_82 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_81;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_83 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_82;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_84 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_83;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_85 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_84;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_86 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_85;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_87 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_86;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_88 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_87;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_89 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_88;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_90 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_89;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_91 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_90;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_92 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_91;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_93 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_92;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_94 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_93;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_95 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_94;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_96 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_95;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_97 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_96;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_98 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_97;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_99 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_98;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_100 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_99;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_101 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_100;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_102 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_101;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_103 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_102;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_104 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_103;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_105 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_104;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_106 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_105;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_107 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_106;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_108 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_107;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_109 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_108;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_110 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_109;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_111 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_110;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_112 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_111;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_113 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_112;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_114 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_113;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_115 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_114;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_116 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_115;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_117 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_116;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_118 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_117;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_119 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_118;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_120 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_119;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_121 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_120;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_122 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_121;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_123 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_122;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_124 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_123;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_125 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_124;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_126 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_125;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_127 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_126;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_128 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_127;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_129 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_128;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_130 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_129;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_131 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_130;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_132 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_131;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_133 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_132;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_134 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_133;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_135 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_134;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_136 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_135;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_137 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_136;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_138 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_137;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_139 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_138;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_140 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_139;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_141 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_140;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_142 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_141;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_143 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_142;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_144 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_143;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_145 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_144;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_146 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_145;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_147 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_146;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_148 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_147;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_149 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_148;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_150 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_149;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_151 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_150;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_152 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_151;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_153 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_152;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_154 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_153;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_155 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_154;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_156 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_155;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_157 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_156;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_158 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_157;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_159 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_158;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_160 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_159;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_161 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_160;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_162 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_161;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_163 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_162;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_164 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_163;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_165 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_164;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_166 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_165;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_167 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_166;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_168 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_167;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_169 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_168;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_170 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_169;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_171 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_170;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_172 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_171;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_173 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_172;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_174 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_173;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_175 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_174;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_176 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_175;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_177 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_176;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_178 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_177;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_179 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_178;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_180 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_179;
      dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_181 <= dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11_stage_180;
      bright_gauss_blur_1_update_0_stage_21 <= bright_gauss_blur_1_update_0;
      bright_gauss_blur_1_update_0_stage_22 <= bright_gauss_blur_1_update_0_stage_21;
      bright_gauss_blur_1_update_0_stage_23 <= bright_gauss_blur_1_update_0_stage_22;
      bright_gauss_blur_1_update_0_stage_24 <= bright_gauss_blur_1_update_0_stage_23;
      bright_gauss_blur_1_update_0_stage_25 <= bright_gauss_blur_1_update_0_stage_24;
      bright_gauss_blur_1_update_0_stage_26 <= bright_gauss_blur_1_update_0_stage_25;
      bright_gauss_blur_1_update_0_stage_27 <= bright_gauss_blur_1_update_0_stage_26;
      bright_gauss_blur_1_update_0_stage_28 <= bright_gauss_blur_1_update_0_stage_27;
      bright_gauss_blur_1_update_0_stage_29 <= bright_gauss_blur_1_update_0_stage_28;
      bright_gauss_blur_1_update_0_stage_30 <= bright_gauss_blur_1_update_0_stage_29;
      bright_gauss_blur_1_update_0_stage_31 <= bright_gauss_blur_1_update_0_stage_30;
      bright_gauss_blur_1_update_0_stage_32 <= bright_gauss_blur_1_update_0_stage_31;
      bright_gauss_blur_1_update_0_stage_33 <= bright_gauss_blur_1_update_0_stage_32;
      bright_gauss_blur_1_update_0_stage_34 <= bright_gauss_blur_1_update_0_stage_33;
      bright_gauss_blur_1_update_0_stage_35 <= bright_gauss_blur_1_update_0_stage_34;
      bright_gauss_blur_1_update_0_stage_36 <= bright_gauss_blur_1_update_0_stage_35;
      bright_gauss_blur_1_update_0_stage_37 <= bright_gauss_blur_1_update_0_stage_36;
      bright_gauss_blur_1_update_0_stage_38 <= bright_gauss_blur_1_update_0_stage_37;
      bright_gauss_blur_1_update_0_stage_39 <= bright_gauss_blur_1_update_0_stage_38;
      bright_gauss_blur_1_update_0_stage_40 <= bright_gauss_blur_1_update_0_stage_39;
      bright_gauss_blur_1_update_0_stage_41 <= bright_gauss_blur_1_update_0_stage_40;
      bright_gauss_blur_1_update_0_stage_42 <= bright_gauss_blur_1_update_0_stage_41;
      bright_gauss_blur_1_update_0_stage_43 <= bright_gauss_blur_1_update_0_stage_42;
      bright_gauss_blur_1_update_0_stage_44 <= bright_gauss_blur_1_update_0_stage_43;
      bright_gauss_blur_1_update_0_stage_45 <= bright_gauss_blur_1_update_0_stage_44;
      bright_gauss_blur_1_update_0_stage_46 <= bright_gauss_blur_1_update_0_stage_45;
      bright_gauss_blur_1_update_0_stage_47 <= bright_gauss_blur_1_update_0_stage_46;
      bright_gauss_blur_1_update_0_stage_48 <= bright_gauss_blur_1_update_0_stage_47;
      bright_gauss_blur_1_update_0_stage_49 <= bright_gauss_blur_1_update_0_stage_48;
      bright_gauss_blur_1_update_0_stage_50 <= bright_gauss_blur_1_update_0_stage_49;
      bright_gauss_blur_1_update_0_stage_51 <= bright_gauss_blur_1_update_0_stage_50;
      bright_gauss_blur_1_update_0_stage_52 <= bright_gauss_blur_1_update_0_stage_51;
      bright_gauss_blur_1_update_0_stage_53 <= bright_gauss_blur_1_update_0_stage_52;
      bright_gauss_blur_1_update_0_stage_54 <= bright_gauss_blur_1_update_0_stage_53;
      bright_gauss_blur_1_update_0_stage_55 <= bright_gauss_blur_1_update_0_stage_54;
      bright_gauss_blur_1_update_0_stage_56 <= bright_gauss_blur_1_update_0_stage_55;
      bright_gauss_blur_1_update_0_stage_57 <= bright_gauss_blur_1_update_0_stage_56;
      bright_gauss_blur_1_update_0_stage_58 <= bright_gauss_blur_1_update_0_stage_57;
      bright_gauss_blur_1_update_0_stage_59 <= bright_gauss_blur_1_update_0_stage_58;
      bright_gauss_blur_1_update_0_stage_60 <= bright_gauss_blur_1_update_0_stage_59;
      bright_gauss_blur_1_update_0_stage_61 <= bright_gauss_blur_1_update_0_stage_60;
      bright_gauss_blur_1_update_0_stage_62 <= bright_gauss_blur_1_update_0_stage_61;
      bright_gauss_blur_1_update_0_stage_63 <= bright_gauss_blur_1_update_0_stage_62;
      bright_gauss_blur_1_update_0_stage_64 <= bright_gauss_blur_1_update_0_stage_63;
      bright_gauss_blur_1_update_0_stage_65 <= bright_gauss_blur_1_update_0_stage_64;
      bright_gauss_blur_1_update_0_stage_66 <= bright_gauss_blur_1_update_0_stage_65;
      bright_gauss_blur_1_update_0_stage_67 <= bright_gauss_blur_1_update_0_stage_66;
      bright_gauss_blur_1_update_0_stage_68 <= bright_gauss_blur_1_update_0_stage_67;
      bright_gauss_blur_1_update_0_stage_69 <= bright_gauss_blur_1_update_0_stage_68;
      bright_gauss_blur_1_update_0_stage_70 <= bright_gauss_blur_1_update_0_stage_69;
      bright_gauss_blur_1_update_0_stage_71 <= bright_gauss_blur_1_update_0_stage_70;
      bright_gauss_blur_1_update_0_stage_72 <= bright_gauss_blur_1_update_0_stage_71;
      bright_gauss_blur_1_update_0_stage_73 <= bright_gauss_blur_1_update_0_stage_72;
      bright_gauss_blur_1_update_0_stage_74 <= bright_gauss_blur_1_update_0_stage_73;
      bright_gauss_blur_1_update_0_stage_75 <= bright_gauss_blur_1_update_0_stage_74;
      bright_gauss_blur_1_update_0_stage_76 <= bright_gauss_blur_1_update_0_stage_75;
      bright_gauss_blur_1_update_0_stage_77 <= bright_gauss_blur_1_update_0_stage_76;
      bright_gauss_blur_1_update_0_stage_78 <= bright_gauss_blur_1_update_0_stage_77;
      bright_gauss_blur_1_update_0_stage_79 <= bright_gauss_blur_1_update_0_stage_78;
      bright_gauss_blur_1_update_0_stage_80 <= bright_gauss_blur_1_update_0_stage_79;
      bright_gauss_blur_1_update_0_stage_81 <= bright_gauss_blur_1_update_0_stage_80;
      bright_gauss_blur_1_update_0_stage_82 <= bright_gauss_blur_1_update_0_stage_81;
      bright_gauss_blur_1_update_0_stage_83 <= bright_gauss_blur_1_update_0_stage_82;
      bright_gauss_blur_1_update_0_stage_84 <= bright_gauss_blur_1_update_0_stage_83;
      bright_gauss_blur_1_update_0_stage_85 <= bright_gauss_blur_1_update_0_stage_84;
      bright_gauss_blur_1_update_0_stage_86 <= bright_gauss_blur_1_update_0_stage_85;
      bright_gauss_blur_1_update_0_stage_87 <= bright_gauss_blur_1_update_0_stage_86;
      bright_gauss_blur_1_update_0_stage_88 <= bright_gauss_blur_1_update_0_stage_87;
      bright_gauss_blur_1_update_0_stage_89 <= bright_gauss_blur_1_update_0_stage_88;
      bright_gauss_blur_1_update_0_stage_90 <= bright_gauss_blur_1_update_0_stage_89;
      bright_gauss_blur_1_update_0_stage_91 <= bright_gauss_blur_1_update_0_stage_90;
      bright_gauss_blur_1_update_0_stage_92 <= bright_gauss_blur_1_update_0_stage_91;
      bright_gauss_blur_1_update_0_stage_93 <= bright_gauss_blur_1_update_0_stage_92;
      bright_gauss_blur_1_update_0_stage_94 <= bright_gauss_blur_1_update_0_stage_93;
      bright_gauss_blur_1_update_0_stage_95 <= bright_gauss_blur_1_update_0_stage_94;
      bright_gauss_blur_1_update_0_stage_96 <= bright_gauss_blur_1_update_0_stage_95;
      bright_gauss_blur_1_update_0_stage_97 <= bright_gauss_blur_1_update_0_stage_96;
      bright_gauss_blur_1_update_0_stage_98 <= bright_gauss_blur_1_update_0_stage_97;
      bright_gauss_blur_1_update_0_stage_99 <= bright_gauss_blur_1_update_0_stage_98;
      bright_gauss_blur_1_update_0_stage_100 <= bright_gauss_blur_1_update_0_stage_99;
      bright_gauss_blur_1_update_0_stage_101 <= bright_gauss_blur_1_update_0_stage_100;
      bright_gauss_blur_1_update_0_stage_102 <= bright_gauss_blur_1_update_0_stage_101;
      bright_gauss_blur_1_update_0_stage_103 <= bright_gauss_blur_1_update_0_stage_102;
      bright_gauss_blur_1_update_0_stage_104 <= bright_gauss_blur_1_update_0_stage_103;
      bright_gauss_blur_1_update_0_stage_105 <= bright_gauss_blur_1_update_0_stage_104;
      bright_gauss_blur_1_update_0_stage_106 <= bright_gauss_blur_1_update_0_stage_105;
      bright_gauss_blur_1_update_0_stage_107 <= bright_gauss_blur_1_update_0_stage_106;
      bright_gauss_blur_1_update_0_stage_108 <= bright_gauss_blur_1_update_0_stage_107;
      bright_gauss_blur_1_update_0_stage_109 <= bright_gauss_blur_1_update_0_stage_108;
      bright_gauss_blur_1_update_0_stage_110 <= bright_gauss_blur_1_update_0_stage_109;
      bright_gauss_blur_1_update_0_stage_111 <= bright_gauss_blur_1_update_0_stage_110;
      bright_gauss_blur_1_update_0_stage_112 <= bright_gauss_blur_1_update_0_stage_111;
      bright_gauss_blur_1_update_0_stage_113 <= bright_gauss_blur_1_update_0_stage_112;
      bright_gauss_blur_1_update_0_stage_114 <= bright_gauss_blur_1_update_0_stage_113;
      bright_gauss_blur_1_update_0_stage_115 <= bright_gauss_blur_1_update_0_stage_114;
      bright_gauss_blur_1_update_0_stage_116 <= bright_gauss_blur_1_update_0_stage_115;
      bright_gauss_blur_1_update_0_stage_117 <= bright_gauss_blur_1_update_0_stage_116;
      bright_gauss_blur_1_update_0_stage_118 <= bright_gauss_blur_1_update_0_stage_117;
      bright_gauss_blur_1_update_0_stage_119 <= bright_gauss_blur_1_update_0_stage_118;
      bright_gauss_blur_1_update_0_stage_120 <= bright_gauss_blur_1_update_0_stage_119;
      bright_gauss_blur_1_update_0_stage_121 <= bright_gauss_blur_1_update_0_stage_120;
      bright_gauss_blur_1_update_0_stage_122 <= bright_gauss_blur_1_update_0_stage_121;
      bright_gauss_blur_1_update_0_stage_123 <= bright_gauss_blur_1_update_0_stage_122;
      bright_gauss_blur_1_update_0_stage_124 <= bright_gauss_blur_1_update_0_stage_123;
      bright_gauss_blur_1_update_0_stage_125 <= bright_gauss_blur_1_update_0_stage_124;
      bright_gauss_blur_1_update_0_stage_126 <= bright_gauss_blur_1_update_0_stage_125;
      bright_gauss_blur_1_update_0_stage_127 <= bright_gauss_blur_1_update_0_stage_126;
      bright_gauss_blur_1_update_0_stage_128 <= bright_gauss_blur_1_update_0_stage_127;
      bright_gauss_blur_1_update_0_stage_129 <= bright_gauss_blur_1_update_0_stage_128;
      bright_gauss_blur_1_update_0_stage_130 <= bright_gauss_blur_1_update_0_stage_129;
      bright_gauss_blur_1_update_0_stage_131 <= bright_gauss_blur_1_update_0_stage_130;
      bright_gauss_blur_1_update_0_stage_132 <= bright_gauss_blur_1_update_0_stage_131;
      bright_gauss_blur_1_update_0_stage_133 <= bright_gauss_blur_1_update_0_stage_132;
      bright_gauss_blur_1_update_0_stage_134 <= bright_gauss_blur_1_update_0_stage_133;
      bright_gauss_blur_1_update_0_stage_135 <= bright_gauss_blur_1_update_0_stage_134;
      bright_gauss_blur_1_update_0_stage_136 <= bright_gauss_blur_1_update_0_stage_135;
      bright_gauss_blur_1_update_0_stage_137 <= bright_gauss_blur_1_update_0_stage_136;
      bright_gauss_blur_1_update_0_stage_138 <= bright_gauss_blur_1_update_0_stage_137;
      bright_gauss_blur_1_update_0_stage_139 <= bright_gauss_blur_1_update_0_stage_138;
      bright_gauss_blur_1_update_0_stage_140 <= bright_gauss_blur_1_update_0_stage_139;
      bright_gauss_blur_1_update_0_stage_141 <= bright_gauss_blur_1_update_0_stage_140;
      bright_gauss_blur_1_update_0_stage_142 <= bright_gauss_blur_1_update_0_stage_141;
      bright_gauss_blur_1_update_0_stage_143 <= bright_gauss_blur_1_update_0_stage_142;
      bright_gauss_blur_1_update_0_stage_144 <= bright_gauss_blur_1_update_0_stage_143;
      bright_gauss_blur_1_update_0_stage_145 <= bright_gauss_blur_1_update_0_stage_144;
      bright_gauss_blur_1_update_0_stage_146 <= bright_gauss_blur_1_update_0_stage_145;
      bright_gauss_blur_1_update_0_stage_147 <= bright_gauss_blur_1_update_0_stage_146;
      bright_gauss_blur_1_update_0_stage_148 <= bright_gauss_blur_1_update_0_stage_147;
      bright_gauss_blur_1_update_0_stage_149 <= bright_gauss_blur_1_update_0_stage_148;
      bright_gauss_blur_1_update_0_stage_150 <= bright_gauss_blur_1_update_0_stage_149;
      bright_gauss_blur_1_update_0_stage_151 <= bright_gauss_blur_1_update_0_stage_150;
      bright_gauss_blur_1_update_0_stage_152 <= bright_gauss_blur_1_update_0_stage_151;
      bright_gauss_blur_1_update_0_stage_153 <= bright_gauss_blur_1_update_0_stage_152;
      bright_gauss_blur_1_update_0_stage_154 <= bright_gauss_blur_1_update_0_stage_153;
      bright_gauss_blur_1_update_0_stage_155 <= bright_gauss_blur_1_update_0_stage_154;
      bright_gauss_blur_1_update_0_stage_156 <= bright_gauss_blur_1_update_0_stage_155;
      bright_gauss_blur_1_update_0_stage_157 <= bright_gauss_blur_1_update_0_stage_156;
      bright_gauss_blur_1_update_0_stage_158 <= bright_gauss_blur_1_update_0_stage_157;
      bright_gauss_blur_1_update_0_stage_159 <= bright_gauss_blur_1_update_0_stage_158;
      bright_gauss_blur_1_update_0_stage_160 <= bright_gauss_blur_1_update_0_stage_159;
      bright_gauss_blur_1_update_0_stage_161 <= bright_gauss_blur_1_update_0_stage_160;
      bright_gauss_blur_1_update_0_stage_162 <= bright_gauss_blur_1_update_0_stage_161;
      bright_gauss_blur_1_update_0_stage_163 <= bright_gauss_blur_1_update_0_stage_162;
      bright_gauss_blur_1_update_0_stage_164 <= bright_gauss_blur_1_update_0_stage_163;
      bright_gauss_blur_1_update_0_stage_165 <= bright_gauss_blur_1_update_0_stage_164;
      bright_gauss_blur_1_update_0_stage_166 <= bright_gauss_blur_1_update_0_stage_165;
      bright_gauss_blur_1_update_0_stage_167 <= bright_gauss_blur_1_update_0_stage_166;
      bright_gauss_blur_1_update_0_stage_168 <= bright_gauss_blur_1_update_0_stage_167;
      bright_gauss_blur_1_update_0_stage_169 <= bright_gauss_blur_1_update_0_stage_168;
      bright_gauss_blur_1_update_0_stage_170 <= bright_gauss_blur_1_update_0_stage_169;
      bright_gauss_blur_1_update_0_stage_171 <= bright_gauss_blur_1_update_0_stage_170;
      bright_gauss_blur_1_update_0_stage_172 <= bright_gauss_blur_1_update_0_stage_171;
      bright_gauss_blur_1_update_0_stage_173 <= bright_gauss_blur_1_update_0_stage_172;
      bright_gauss_blur_1_update_0_stage_174 <= bright_gauss_blur_1_update_0_stage_173;
      bright_gauss_blur_1_update_0_stage_175 <= bright_gauss_blur_1_update_0_stage_174;
      bright_gauss_blur_1_update_0_stage_176 <= bright_gauss_blur_1_update_0_stage_175;
      bright_gauss_blur_1_update_0_stage_177 <= bright_gauss_blur_1_update_0_stage_176;
      bright_gauss_blur_1_update_0_stage_178 <= bright_gauss_blur_1_update_0_stage_177;
      bright_gauss_blur_1_update_0_stage_179 <= bright_gauss_blur_1_update_0_stage_178;
      bright_gauss_blur_1_update_0_stage_180 <= bright_gauss_blur_1_update_0_stage_179;
      bright_gauss_blur_1_update_0_stage_181 <= bright_gauss_blur_1_update_0_stage_180;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_20 <= bright_bright_gauss_blur_1_update_0_read_read_12;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_21 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_20;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_22 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_21;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_23 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_22;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_24 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_23;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_25 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_24;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_26 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_25;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_27 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_26;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_28 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_27;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_29 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_28;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_30 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_29;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_31 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_30;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_32 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_31;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_33 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_32;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_34 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_33;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_35 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_34;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_36 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_35;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_37 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_36;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_38 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_37;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_39 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_38;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_40 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_39;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_41 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_40;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_42 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_41;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_43 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_42;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_44 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_43;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_45 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_44;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_46 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_45;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_47 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_46;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_48 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_47;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_49 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_48;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_50 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_49;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_51 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_50;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_52 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_51;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_53 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_52;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_54 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_53;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_55 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_54;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_56 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_55;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_57 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_56;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_58 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_57;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_59 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_58;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_60 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_59;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_61 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_60;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_62 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_61;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_63 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_62;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_64 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_63;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_65 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_64;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_66 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_65;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_67 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_66;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_68 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_67;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_69 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_68;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_70 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_69;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_71 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_70;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_72 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_71;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_73 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_72;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_74 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_73;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_75 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_74;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_76 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_75;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_77 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_76;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_78 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_77;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_79 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_78;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_80 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_79;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_81 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_80;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_82 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_81;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_83 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_82;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_84 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_83;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_85 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_84;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_86 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_85;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_87 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_86;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_88 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_87;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_89 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_88;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_90 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_89;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_91 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_90;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_92 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_91;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_93 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_92;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_94 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_93;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_95 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_94;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_96 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_95;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_97 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_96;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_98 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_97;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_99 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_98;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_100 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_99;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_101 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_100;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_102 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_101;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_103 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_102;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_104 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_103;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_105 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_104;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_106 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_105;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_107 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_106;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_108 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_107;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_109 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_108;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_110 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_109;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_111 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_110;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_112 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_111;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_113 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_112;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_114 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_113;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_115 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_114;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_116 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_115;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_117 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_116;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_118 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_117;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_119 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_118;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_120 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_119;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_121 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_120;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_122 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_121;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_123 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_122;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_124 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_123;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_125 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_124;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_126 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_125;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_127 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_126;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_128 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_127;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_129 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_128;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_130 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_129;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_131 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_130;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_132 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_131;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_133 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_132;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_134 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_133;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_135 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_134;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_136 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_135;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_137 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_136;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_138 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_137;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_139 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_138;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_140 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_139;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_141 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_140;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_142 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_141;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_143 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_142;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_144 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_143;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_145 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_144;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_146 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_145;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_147 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_146;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_148 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_147;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_149 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_148;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_150 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_149;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_151 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_150;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_152 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_151;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_153 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_152;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_154 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_153;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_155 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_154;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_156 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_155;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_157 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_156;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_158 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_157;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_159 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_158;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_160 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_159;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_161 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_160;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_162 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_161;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_163 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_162;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_164 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_163;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_165 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_164;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_166 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_165;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_167 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_166;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_168 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_167;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_169 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_168;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_170 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_169;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_171 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_170;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_172 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_171;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_173 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_172;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_174 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_173;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_175 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_174;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_176 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_175;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_177 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_176;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_178 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_177;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_179 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_178;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_180 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_179;
      bright_bright_gauss_blur_1_update_0_read_read_12_stage_181 <= bright_bright_gauss_blur_1_update_0_read_read_12_stage_180;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_22 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_23 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_22;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_24 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_23;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_25 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_24;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_26 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_25;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_27 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_26;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_28 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_27;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_29 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_28;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_30 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_29;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_31 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_30;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_32 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_31;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_33 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_32;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_34 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_33;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_35 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_34;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_36 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_35;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_37 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_36;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_38 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_37;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_39 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_38;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_40 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_39;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_41 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_40;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_42 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_41;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_43 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_42;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_44 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_43;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_45 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_44;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_46 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_45;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_47 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_46;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_48 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_47;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_49 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_48;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_50 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_49;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_51 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_50;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_52 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_51;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_53 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_52;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_54 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_53;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_55 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_54;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_56 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_55;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_57 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_56;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_58 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_57;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_59 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_58;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_60 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_59;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_61 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_60;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_62 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_61;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_63 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_62;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_64 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_63;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_65 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_64;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_66 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_65;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_67 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_66;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_68 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_67;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_69 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_68;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_70 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_69;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_71 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_70;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_72 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_71;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_73 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_72;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_74 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_73;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_75 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_74;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_76 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_75;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_77 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_76;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_78 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_77;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_79 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_78;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_80 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_79;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_81 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_80;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_82 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_81;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_83 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_82;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_84 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_83;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_85 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_84;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_86 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_85;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_87 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_86;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_88 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_87;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_89 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_88;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_90 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_89;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_91 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_90;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_92 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_91;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_93 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_92;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_94 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_93;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_95 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_94;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_96 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_95;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_97 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_96;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_98 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_97;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_99 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_98;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_100 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_99;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_101 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_100;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_102 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_101;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_103 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_102;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_104 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_103;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_105 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_104;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_106 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_105;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_107 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_106;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_108 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_107;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_109 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_108;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_110 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_109;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_111 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_110;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_112 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_111;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_113 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_112;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_114 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_113;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_115 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_114;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_116 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_115;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_117 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_116;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_118 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_117;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_119 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_118;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_120 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_119;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_121 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_120;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_122 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_121;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_123 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_122;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_124 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_123;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_125 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_124;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_126 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_125;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_127 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_126;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_128 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_127;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_129 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_128;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_130 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_129;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_131 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_130;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_132 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_131;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_133 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_132;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_134 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_133;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_135 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_134;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_136 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_135;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_137 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_136;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_138 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_137;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_139 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_138;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_140 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_139;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_141 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_140;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_142 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_141;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_143 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_142;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_144 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_143;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_145 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_144;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_146 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_145;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_147 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_146;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_148 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_147;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_149 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_148;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_150 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_149;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_151 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_150;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_152 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_151;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_153 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_152;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_154 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_153;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_155 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_154;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_156 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_155;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_157 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_156;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_158 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_157;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_159 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_158;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_160 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_159;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_161 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_160;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_162 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_161;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_163 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_162;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_164 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_163;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_165 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_164;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_166 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_165;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_167 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_166;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_168 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_167;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_169 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_168;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_170 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_169;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_171 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_170;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_172 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_171;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_173 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_172;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_174 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_173;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_175 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_174;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_176 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_175;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_177 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_176;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_178 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_177;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_179 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_178;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_180 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_179;
      bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_181 <= bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13_stage_180;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_61 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_62 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_61;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_63 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_62;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_64 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_63;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_65 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_64;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_66 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_65;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_67 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_66;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_68 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_67;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_69 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_68;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_70 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_69;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_71 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_70;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_72 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_71;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_73 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_72;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_74 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_73;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_75 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_74;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_76 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_75;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_77 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_76;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_78 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_77;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_79 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_78;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_80 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_79;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_81 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_80;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_82 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_81;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_83 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_82;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_84 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_83;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_85 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_84;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_86 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_85;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_87 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_86;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_88 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_87;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_89 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_88;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_90 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_89;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_91 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_90;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_92 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_91;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_93 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_92;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_94 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_93;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_95 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_94;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_96 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_95;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_97 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_96;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_98 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_97;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_99 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_98;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_100 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_99;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_101 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_100;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_102 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_101;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_103 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_102;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_104 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_103;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_105 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_104;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_106 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_105;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_107 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_106;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_108 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_107;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_109 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_108;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_110 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_109;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_111 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_110;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_112 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_111;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_113 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_112;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_114 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_113;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_115 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_114;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_116 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_115;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_117 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_116;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_118 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_117;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_119 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_118;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_120 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_119;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_121 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_120;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_122 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_121;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_123 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_122;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_124 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_123;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_125 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_124;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_126 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_125;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_127 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_126;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_128 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_127;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_129 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_128;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_130 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_129;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_131 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_130;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_132 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_131;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_133 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_132;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_134 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_133;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_135 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_134;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_136 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_135;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_137 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_136;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_138 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_137;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_139 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_138;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_140 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_139;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_141 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_140;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_142 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_141;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_143 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_142;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_144 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_143;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_145 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_144;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_146 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_145;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_147 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_146;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_148 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_147;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_149 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_148;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_150 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_149;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_151 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_150;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_152 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_151;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_153 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_152;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_154 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_153;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_155 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_154;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_156 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_155;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_157 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_156;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_158 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_157;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_159 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_158;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_160 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_159;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_161 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_160;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_162 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_161;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_163 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_162;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_164 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_163;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_165 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_164;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_166 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_165;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_167 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_166;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_168 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_167;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_169 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_168;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_170 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_169;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_171 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_170;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_172 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_171;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_173 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_172;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_174 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_173;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_175 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_174;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_176 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_175;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_177 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_176;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_178 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_177;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_179 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_178;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_180 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_179;
      bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_181 <= bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40_stage_180;
      bright_laplace_us_1_update_0_stage_62 <= bright_laplace_us_1_update_0;
      bright_laplace_us_1_update_0_stage_63 <= bright_laplace_us_1_update_0_stage_62;
      bright_laplace_us_1_update_0_stage_64 <= bright_laplace_us_1_update_0_stage_63;
      bright_laplace_us_1_update_0_stage_65 <= bright_laplace_us_1_update_0_stage_64;
      bright_laplace_us_1_update_0_stage_66 <= bright_laplace_us_1_update_0_stage_65;
      bright_laplace_us_1_update_0_stage_67 <= bright_laplace_us_1_update_0_stage_66;
      bright_laplace_us_1_update_0_stage_68 <= bright_laplace_us_1_update_0_stage_67;
      bright_laplace_us_1_update_0_stage_69 <= bright_laplace_us_1_update_0_stage_68;
      bright_laplace_us_1_update_0_stage_70 <= bright_laplace_us_1_update_0_stage_69;
      bright_laplace_us_1_update_0_stage_71 <= bright_laplace_us_1_update_0_stage_70;
      bright_laplace_us_1_update_0_stage_72 <= bright_laplace_us_1_update_0_stage_71;
      bright_laplace_us_1_update_0_stage_73 <= bright_laplace_us_1_update_0_stage_72;
      bright_laplace_us_1_update_0_stage_74 <= bright_laplace_us_1_update_0_stage_73;
      bright_laplace_us_1_update_0_stage_75 <= bright_laplace_us_1_update_0_stage_74;
      bright_laplace_us_1_update_0_stage_76 <= bright_laplace_us_1_update_0_stage_75;
      bright_laplace_us_1_update_0_stage_77 <= bright_laplace_us_1_update_0_stage_76;
      bright_laplace_us_1_update_0_stage_78 <= bright_laplace_us_1_update_0_stage_77;
      bright_laplace_us_1_update_0_stage_79 <= bright_laplace_us_1_update_0_stage_78;
      bright_laplace_us_1_update_0_stage_80 <= bright_laplace_us_1_update_0_stage_79;
      bright_laplace_us_1_update_0_stage_81 <= bright_laplace_us_1_update_0_stage_80;
      bright_laplace_us_1_update_0_stage_82 <= bright_laplace_us_1_update_0_stage_81;
      bright_laplace_us_1_update_0_stage_83 <= bright_laplace_us_1_update_0_stage_82;
      bright_laplace_us_1_update_0_stage_84 <= bright_laplace_us_1_update_0_stage_83;
      bright_laplace_us_1_update_0_stage_85 <= bright_laplace_us_1_update_0_stage_84;
      bright_laplace_us_1_update_0_stage_86 <= bright_laplace_us_1_update_0_stage_85;
      bright_laplace_us_1_update_0_stage_87 <= bright_laplace_us_1_update_0_stage_86;
      bright_laplace_us_1_update_0_stage_88 <= bright_laplace_us_1_update_0_stage_87;
      bright_laplace_us_1_update_0_stage_89 <= bright_laplace_us_1_update_0_stage_88;
      bright_laplace_us_1_update_0_stage_90 <= bright_laplace_us_1_update_0_stage_89;
      bright_laplace_us_1_update_0_stage_91 <= bright_laplace_us_1_update_0_stage_90;
      bright_laplace_us_1_update_0_stage_92 <= bright_laplace_us_1_update_0_stage_91;
      bright_laplace_us_1_update_0_stage_93 <= bright_laplace_us_1_update_0_stage_92;
      bright_laplace_us_1_update_0_stage_94 <= bright_laplace_us_1_update_0_stage_93;
      bright_laplace_us_1_update_0_stage_95 <= bright_laplace_us_1_update_0_stage_94;
      bright_laplace_us_1_update_0_stage_96 <= bright_laplace_us_1_update_0_stage_95;
      bright_laplace_us_1_update_0_stage_97 <= bright_laplace_us_1_update_0_stage_96;
      bright_laplace_us_1_update_0_stage_98 <= bright_laplace_us_1_update_0_stage_97;
      bright_laplace_us_1_update_0_stage_99 <= bright_laplace_us_1_update_0_stage_98;
      bright_laplace_us_1_update_0_stage_100 <= bright_laplace_us_1_update_0_stage_99;
      bright_laplace_us_1_update_0_stage_101 <= bright_laplace_us_1_update_0_stage_100;
      bright_laplace_us_1_update_0_stage_102 <= bright_laplace_us_1_update_0_stage_101;
      bright_laplace_us_1_update_0_stage_103 <= bright_laplace_us_1_update_0_stage_102;
      bright_laplace_us_1_update_0_stage_104 <= bright_laplace_us_1_update_0_stage_103;
      bright_laplace_us_1_update_0_stage_105 <= bright_laplace_us_1_update_0_stage_104;
      bright_laplace_us_1_update_0_stage_106 <= bright_laplace_us_1_update_0_stage_105;
      bright_laplace_us_1_update_0_stage_107 <= bright_laplace_us_1_update_0_stage_106;
      bright_laplace_us_1_update_0_stage_108 <= bright_laplace_us_1_update_0_stage_107;
      bright_laplace_us_1_update_0_stage_109 <= bright_laplace_us_1_update_0_stage_108;
      bright_laplace_us_1_update_0_stage_110 <= bright_laplace_us_1_update_0_stage_109;
      bright_laplace_us_1_update_0_stage_111 <= bright_laplace_us_1_update_0_stage_110;
      bright_laplace_us_1_update_0_stage_112 <= bright_laplace_us_1_update_0_stage_111;
      bright_laplace_us_1_update_0_stage_113 <= bright_laplace_us_1_update_0_stage_112;
      bright_laplace_us_1_update_0_stage_114 <= bright_laplace_us_1_update_0_stage_113;
      bright_laplace_us_1_update_0_stage_115 <= bright_laplace_us_1_update_0_stage_114;
      bright_laplace_us_1_update_0_stage_116 <= bright_laplace_us_1_update_0_stage_115;
      bright_laplace_us_1_update_0_stage_117 <= bright_laplace_us_1_update_0_stage_116;
      bright_laplace_us_1_update_0_stage_118 <= bright_laplace_us_1_update_0_stage_117;
      bright_laplace_us_1_update_0_stage_119 <= bright_laplace_us_1_update_0_stage_118;
      bright_laplace_us_1_update_0_stage_120 <= bright_laplace_us_1_update_0_stage_119;
      bright_laplace_us_1_update_0_stage_121 <= bright_laplace_us_1_update_0_stage_120;
      bright_laplace_us_1_update_0_stage_122 <= bright_laplace_us_1_update_0_stage_121;
      bright_laplace_us_1_update_0_stage_123 <= bright_laplace_us_1_update_0_stage_122;
      bright_laplace_us_1_update_0_stage_124 <= bright_laplace_us_1_update_0_stage_123;
      bright_laplace_us_1_update_0_stage_125 <= bright_laplace_us_1_update_0_stage_124;
      bright_laplace_us_1_update_0_stage_126 <= bright_laplace_us_1_update_0_stage_125;
      bright_laplace_us_1_update_0_stage_127 <= bright_laplace_us_1_update_0_stage_126;
      bright_laplace_us_1_update_0_stage_128 <= bright_laplace_us_1_update_0_stage_127;
      bright_laplace_us_1_update_0_stage_129 <= bright_laplace_us_1_update_0_stage_128;
      bright_laplace_us_1_update_0_stage_130 <= bright_laplace_us_1_update_0_stage_129;
      bright_laplace_us_1_update_0_stage_131 <= bright_laplace_us_1_update_0_stage_130;
      bright_laplace_us_1_update_0_stage_132 <= bright_laplace_us_1_update_0_stage_131;
      bright_laplace_us_1_update_0_stage_133 <= bright_laplace_us_1_update_0_stage_132;
      bright_laplace_us_1_update_0_stage_134 <= bright_laplace_us_1_update_0_stage_133;
      bright_laplace_us_1_update_0_stage_135 <= bright_laplace_us_1_update_0_stage_134;
      bright_laplace_us_1_update_0_stage_136 <= bright_laplace_us_1_update_0_stage_135;
      bright_laplace_us_1_update_0_stage_137 <= bright_laplace_us_1_update_0_stage_136;
      bright_laplace_us_1_update_0_stage_138 <= bright_laplace_us_1_update_0_stage_137;
      bright_laplace_us_1_update_0_stage_139 <= bright_laplace_us_1_update_0_stage_138;
      bright_laplace_us_1_update_0_stage_140 <= bright_laplace_us_1_update_0_stage_139;
      bright_laplace_us_1_update_0_stage_141 <= bright_laplace_us_1_update_0_stage_140;
      bright_laplace_us_1_update_0_stage_142 <= bright_laplace_us_1_update_0_stage_141;
      bright_laplace_us_1_update_0_stage_143 <= bright_laplace_us_1_update_0_stage_142;
      bright_laplace_us_1_update_0_stage_144 <= bright_laplace_us_1_update_0_stage_143;
      bright_laplace_us_1_update_0_stage_145 <= bright_laplace_us_1_update_0_stage_144;
      bright_laplace_us_1_update_0_stage_146 <= bright_laplace_us_1_update_0_stage_145;
      bright_laplace_us_1_update_0_stage_147 <= bright_laplace_us_1_update_0_stage_146;
      bright_laplace_us_1_update_0_stage_148 <= bright_laplace_us_1_update_0_stage_147;
      bright_laplace_us_1_update_0_stage_149 <= bright_laplace_us_1_update_0_stage_148;
      bright_laplace_us_1_update_0_stage_150 <= bright_laplace_us_1_update_0_stage_149;
      bright_laplace_us_1_update_0_stage_151 <= bright_laplace_us_1_update_0_stage_150;
      bright_laplace_us_1_update_0_stage_152 <= bright_laplace_us_1_update_0_stage_151;
      bright_laplace_us_1_update_0_stage_153 <= bright_laplace_us_1_update_0_stage_152;
      bright_laplace_us_1_update_0_stage_154 <= bright_laplace_us_1_update_0_stage_153;
      bright_laplace_us_1_update_0_stage_155 <= bright_laplace_us_1_update_0_stage_154;
      bright_laplace_us_1_update_0_stage_156 <= bright_laplace_us_1_update_0_stage_155;
      bright_laplace_us_1_update_0_stage_157 <= bright_laplace_us_1_update_0_stage_156;
      bright_laplace_us_1_update_0_stage_158 <= bright_laplace_us_1_update_0_stage_157;
      bright_laplace_us_1_update_0_stage_159 <= bright_laplace_us_1_update_0_stage_158;
      bright_laplace_us_1_update_0_stage_160 <= bright_laplace_us_1_update_0_stage_159;
      bright_laplace_us_1_update_0_stage_161 <= bright_laplace_us_1_update_0_stage_160;
      bright_laplace_us_1_update_0_stage_162 <= bright_laplace_us_1_update_0_stage_161;
      bright_laplace_us_1_update_0_stage_163 <= bright_laplace_us_1_update_0_stage_162;
      bright_laplace_us_1_update_0_stage_164 <= bright_laplace_us_1_update_0_stage_163;
      bright_laplace_us_1_update_0_stage_165 <= bright_laplace_us_1_update_0_stage_164;
      bright_laplace_us_1_update_0_stage_166 <= bright_laplace_us_1_update_0_stage_165;
      bright_laplace_us_1_update_0_stage_167 <= bright_laplace_us_1_update_0_stage_166;
      bright_laplace_us_1_update_0_stage_168 <= bright_laplace_us_1_update_0_stage_167;
      bright_laplace_us_1_update_0_stage_169 <= bright_laplace_us_1_update_0_stage_168;
      bright_laplace_us_1_update_0_stage_170 <= bright_laplace_us_1_update_0_stage_169;
      bright_laplace_us_1_update_0_stage_171 <= bright_laplace_us_1_update_0_stage_170;
      bright_laplace_us_1_update_0_stage_172 <= bright_laplace_us_1_update_0_stage_171;
      bright_laplace_us_1_update_0_stage_173 <= bright_laplace_us_1_update_0_stage_172;
      bright_laplace_us_1_update_0_stage_174 <= bright_laplace_us_1_update_0_stage_173;
      bright_laplace_us_1_update_0_stage_175 <= bright_laplace_us_1_update_0_stage_174;
      bright_laplace_us_1_update_0_stage_176 <= bright_laplace_us_1_update_0_stage_175;
      bright_laplace_us_1_update_0_stage_177 <= bright_laplace_us_1_update_0_stage_176;
      bright_laplace_us_1_update_0_stage_178 <= bright_laplace_us_1_update_0_stage_177;
      bright_laplace_us_1_update_0_stage_179 <= bright_laplace_us_1_update_0_stage_178;
      bright_laplace_us_1_update_0_stage_180 <= bright_laplace_us_1_update_0_stage_179;
      bright_laplace_us_1_update_0_stage_181 <= bright_laplace_us_1_update_0_stage_180;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_63 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_64 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_63;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_65 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_64;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_66 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_65;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_67 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_66;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_68 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_67;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_69 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_68;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_70 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_69;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_71 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_70;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_72 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_71;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_73 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_72;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_74 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_73;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_75 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_74;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_76 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_75;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_77 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_76;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_78 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_77;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_79 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_78;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_80 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_79;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_81 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_80;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_82 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_81;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_83 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_82;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_84 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_83;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_85 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_84;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_86 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_85;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_87 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_86;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_88 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_87;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_89 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_88;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_90 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_89;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_91 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_90;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_92 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_91;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_93 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_92;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_94 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_93;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_95 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_94;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_96 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_95;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_97 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_96;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_98 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_97;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_99 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_98;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_100 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_99;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_101 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_100;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_102 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_101;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_103 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_102;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_104 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_103;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_105 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_104;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_106 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_105;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_107 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_106;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_108 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_107;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_109 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_108;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_110 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_109;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_111 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_110;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_112 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_111;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_113 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_112;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_114 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_113;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_115 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_114;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_116 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_115;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_117 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_116;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_118 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_117;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_119 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_118;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_120 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_119;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_121 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_120;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_122 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_121;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_123 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_122;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_124 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_123;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_125 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_124;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_126 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_125;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_127 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_126;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_128 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_127;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_129 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_128;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_130 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_129;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_131 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_130;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_132 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_131;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_133 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_132;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_134 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_133;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_135 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_134;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_136 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_135;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_137 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_136;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_138 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_137;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_139 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_138;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_140 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_139;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_141 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_140;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_142 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_141;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_143 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_142;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_144 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_143;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_145 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_144;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_146 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_145;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_147 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_146;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_148 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_147;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_149 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_148;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_150 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_149;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_151 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_150;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_152 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_151;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_153 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_152;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_154 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_153;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_155 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_154;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_156 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_155;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_157 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_156;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_158 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_157;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_159 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_158;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_160 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_159;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_161 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_160;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_162 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_161;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_163 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_162;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_164 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_163;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_165 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_164;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_166 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_165;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_167 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_166;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_168 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_167;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_169 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_168;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_170 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_169;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_171 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_170;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_172 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_171;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_173 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_172;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_174 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_173;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_175 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_174;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_176 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_175;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_177 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_176;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_178 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_177;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_179 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_178;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_180 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_179;
      bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_181 <= bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41_stage_180;
      bright_weights_normed_gauss_blur_1_update_0_stage_83 <= bright_weights_normed_gauss_blur_1_update_0;
      bright_weights_normed_gauss_blur_1_update_0_stage_84 <= bright_weights_normed_gauss_blur_1_update_0_stage_83;
      bright_weights_normed_gauss_blur_1_update_0_stage_85 <= bright_weights_normed_gauss_blur_1_update_0_stage_84;
      bright_weights_normed_gauss_blur_1_update_0_stage_86 <= bright_weights_normed_gauss_blur_1_update_0_stage_85;
      bright_weights_normed_gauss_blur_1_update_0_stage_87 <= bright_weights_normed_gauss_blur_1_update_0_stage_86;
      bright_weights_normed_gauss_blur_1_update_0_stage_88 <= bright_weights_normed_gauss_blur_1_update_0_stage_87;
      bright_weights_normed_gauss_blur_1_update_0_stage_89 <= bright_weights_normed_gauss_blur_1_update_0_stage_88;
      bright_weights_normed_gauss_blur_1_update_0_stage_90 <= bright_weights_normed_gauss_blur_1_update_0_stage_89;
      bright_weights_normed_gauss_blur_1_update_0_stage_91 <= bright_weights_normed_gauss_blur_1_update_0_stage_90;
      bright_weights_normed_gauss_blur_1_update_0_stage_92 <= bright_weights_normed_gauss_blur_1_update_0_stage_91;
      bright_weights_normed_gauss_blur_1_update_0_stage_93 <= bright_weights_normed_gauss_blur_1_update_0_stage_92;
      bright_weights_normed_gauss_blur_1_update_0_stage_94 <= bright_weights_normed_gauss_blur_1_update_0_stage_93;
      bright_weights_normed_gauss_blur_1_update_0_stage_95 <= bright_weights_normed_gauss_blur_1_update_0_stage_94;
      bright_weights_normed_gauss_blur_1_update_0_stage_96 <= bright_weights_normed_gauss_blur_1_update_0_stage_95;
      bright_weights_normed_gauss_blur_1_update_0_stage_97 <= bright_weights_normed_gauss_blur_1_update_0_stage_96;
      bright_weights_normed_gauss_blur_1_update_0_stage_98 <= bright_weights_normed_gauss_blur_1_update_0_stage_97;
      bright_weights_normed_gauss_blur_1_update_0_stage_99 <= bright_weights_normed_gauss_blur_1_update_0_stage_98;
      bright_weights_normed_gauss_blur_1_update_0_stage_100 <= bright_weights_normed_gauss_blur_1_update_0_stage_99;
      bright_weights_normed_gauss_blur_1_update_0_stage_101 <= bright_weights_normed_gauss_blur_1_update_0_stage_100;
      bright_weights_normed_gauss_blur_1_update_0_stage_102 <= bright_weights_normed_gauss_blur_1_update_0_stage_101;
      bright_weights_normed_gauss_blur_1_update_0_stage_103 <= bright_weights_normed_gauss_blur_1_update_0_stage_102;
      bright_weights_normed_gauss_blur_1_update_0_stage_104 <= bright_weights_normed_gauss_blur_1_update_0_stage_103;
      bright_weights_normed_gauss_blur_1_update_0_stage_105 <= bright_weights_normed_gauss_blur_1_update_0_stage_104;
      bright_weights_normed_gauss_blur_1_update_0_stage_106 <= bright_weights_normed_gauss_blur_1_update_0_stage_105;
      bright_weights_normed_gauss_blur_1_update_0_stage_107 <= bright_weights_normed_gauss_blur_1_update_0_stage_106;
      bright_weights_normed_gauss_blur_1_update_0_stage_108 <= bright_weights_normed_gauss_blur_1_update_0_stage_107;
      bright_weights_normed_gauss_blur_1_update_0_stage_109 <= bright_weights_normed_gauss_blur_1_update_0_stage_108;
      bright_weights_normed_gauss_blur_1_update_0_stage_110 <= bright_weights_normed_gauss_blur_1_update_0_stage_109;
      bright_weights_normed_gauss_blur_1_update_0_stage_111 <= bright_weights_normed_gauss_blur_1_update_0_stage_110;
      bright_weights_normed_gauss_blur_1_update_0_stage_112 <= bright_weights_normed_gauss_blur_1_update_0_stage_111;
      bright_weights_normed_gauss_blur_1_update_0_stage_113 <= bright_weights_normed_gauss_blur_1_update_0_stage_112;
      bright_weights_normed_gauss_blur_1_update_0_stage_114 <= bright_weights_normed_gauss_blur_1_update_0_stage_113;
      bright_weights_normed_gauss_blur_1_update_0_stage_115 <= bright_weights_normed_gauss_blur_1_update_0_stage_114;
      bright_weights_normed_gauss_blur_1_update_0_stage_116 <= bright_weights_normed_gauss_blur_1_update_0_stage_115;
      bright_weights_normed_gauss_blur_1_update_0_stage_117 <= bright_weights_normed_gauss_blur_1_update_0_stage_116;
      bright_weights_normed_gauss_blur_1_update_0_stage_118 <= bright_weights_normed_gauss_blur_1_update_0_stage_117;
      bright_weights_normed_gauss_blur_1_update_0_stage_119 <= bright_weights_normed_gauss_blur_1_update_0_stage_118;
      bright_weights_normed_gauss_blur_1_update_0_stage_120 <= bright_weights_normed_gauss_blur_1_update_0_stage_119;
      bright_weights_normed_gauss_blur_1_update_0_stage_121 <= bright_weights_normed_gauss_blur_1_update_0_stage_120;
      bright_weights_normed_gauss_blur_1_update_0_stage_122 <= bright_weights_normed_gauss_blur_1_update_0_stage_121;
      bright_weights_normed_gauss_blur_1_update_0_stage_123 <= bright_weights_normed_gauss_blur_1_update_0_stage_122;
      bright_weights_normed_gauss_blur_1_update_0_stage_124 <= bright_weights_normed_gauss_blur_1_update_0_stage_123;
      bright_weights_normed_gauss_blur_1_update_0_stage_125 <= bright_weights_normed_gauss_blur_1_update_0_stage_124;
      bright_weights_normed_gauss_blur_1_update_0_stage_126 <= bright_weights_normed_gauss_blur_1_update_0_stage_125;
      bright_weights_normed_gauss_blur_1_update_0_stage_127 <= bright_weights_normed_gauss_blur_1_update_0_stage_126;
      bright_weights_normed_gauss_blur_1_update_0_stage_128 <= bright_weights_normed_gauss_blur_1_update_0_stage_127;
      bright_weights_normed_gauss_blur_1_update_0_stage_129 <= bright_weights_normed_gauss_blur_1_update_0_stage_128;
      bright_weights_normed_gauss_blur_1_update_0_stage_130 <= bright_weights_normed_gauss_blur_1_update_0_stage_129;
      bright_weights_normed_gauss_blur_1_update_0_stage_131 <= bright_weights_normed_gauss_blur_1_update_0_stage_130;
      bright_weights_normed_gauss_blur_1_update_0_stage_132 <= bright_weights_normed_gauss_blur_1_update_0_stage_131;
      bright_weights_normed_gauss_blur_1_update_0_stage_133 <= bright_weights_normed_gauss_blur_1_update_0_stage_132;
      bright_weights_normed_gauss_blur_1_update_0_stage_134 <= bright_weights_normed_gauss_blur_1_update_0_stage_133;
      bright_weights_normed_gauss_blur_1_update_0_stage_135 <= bright_weights_normed_gauss_blur_1_update_0_stage_134;
      bright_weights_normed_gauss_blur_1_update_0_stage_136 <= bright_weights_normed_gauss_blur_1_update_0_stage_135;
      bright_weights_normed_gauss_blur_1_update_0_stage_137 <= bright_weights_normed_gauss_blur_1_update_0_stage_136;
      bright_weights_normed_gauss_blur_1_update_0_stage_138 <= bright_weights_normed_gauss_blur_1_update_0_stage_137;
      bright_weights_normed_gauss_blur_1_update_0_stage_139 <= bright_weights_normed_gauss_blur_1_update_0_stage_138;
      bright_weights_normed_gauss_blur_1_update_0_stage_140 <= bright_weights_normed_gauss_blur_1_update_0_stage_139;
      bright_weights_normed_gauss_blur_1_update_0_stage_141 <= bright_weights_normed_gauss_blur_1_update_0_stage_140;
      bright_weights_normed_gauss_blur_1_update_0_stage_142 <= bright_weights_normed_gauss_blur_1_update_0_stage_141;
      bright_weights_normed_gauss_blur_1_update_0_stage_143 <= bright_weights_normed_gauss_blur_1_update_0_stage_142;
      bright_weights_normed_gauss_blur_1_update_0_stage_144 <= bright_weights_normed_gauss_blur_1_update_0_stage_143;
      bright_weights_normed_gauss_blur_1_update_0_stage_145 <= bright_weights_normed_gauss_blur_1_update_0_stage_144;
      bright_weights_normed_gauss_blur_1_update_0_stage_146 <= bright_weights_normed_gauss_blur_1_update_0_stage_145;
      bright_weights_normed_gauss_blur_1_update_0_stage_147 <= bright_weights_normed_gauss_blur_1_update_0_stage_146;
      bright_weights_normed_gauss_blur_1_update_0_stage_148 <= bright_weights_normed_gauss_blur_1_update_0_stage_147;
      bright_weights_normed_gauss_blur_1_update_0_stage_149 <= bright_weights_normed_gauss_blur_1_update_0_stage_148;
      bright_weights_normed_gauss_blur_1_update_0_stage_150 <= bright_weights_normed_gauss_blur_1_update_0_stage_149;
      bright_weights_normed_gauss_blur_1_update_0_stage_151 <= bright_weights_normed_gauss_blur_1_update_0_stage_150;
      bright_weights_normed_gauss_blur_1_update_0_stage_152 <= bright_weights_normed_gauss_blur_1_update_0_stage_151;
      bright_weights_normed_gauss_blur_1_update_0_stage_153 <= bright_weights_normed_gauss_blur_1_update_0_stage_152;
      bright_weights_normed_gauss_blur_1_update_0_stage_154 <= bright_weights_normed_gauss_blur_1_update_0_stage_153;
      bright_weights_normed_gauss_blur_1_update_0_stage_155 <= bright_weights_normed_gauss_blur_1_update_0_stage_154;
      bright_weights_normed_gauss_blur_1_update_0_stage_156 <= bright_weights_normed_gauss_blur_1_update_0_stage_155;
      bright_weights_normed_gauss_blur_1_update_0_stage_157 <= bright_weights_normed_gauss_blur_1_update_0_stage_156;
      bright_weights_normed_gauss_blur_1_update_0_stage_158 <= bright_weights_normed_gauss_blur_1_update_0_stage_157;
      bright_weights_normed_gauss_blur_1_update_0_stage_159 <= bright_weights_normed_gauss_blur_1_update_0_stage_158;
      bright_weights_normed_gauss_blur_1_update_0_stage_160 <= bright_weights_normed_gauss_blur_1_update_0_stage_159;
      bright_weights_normed_gauss_blur_1_update_0_stage_161 <= bright_weights_normed_gauss_blur_1_update_0_stage_160;
      bright_weights_normed_gauss_blur_1_update_0_stage_162 <= bright_weights_normed_gauss_blur_1_update_0_stage_161;
      bright_weights_normed_gauss_blur_1_update_0_stage_163 <= bright_weights_normed_gauss_blur_1_update_0_stage_162;
      bright_weights_normed_gauss_blur_1_update_0_stage_164 <= bright_weights_normed_gauss_blur_1_update_0_stage_163;
      bright_weights_normed_gauss_blur_1_update_0_stage_165 <= bright_weights_normed_gauss_blur_1_update_0_stage_164;
      bright_weights_normed_gauss_blur_1_update_0_stage_166 <= bright_weights_normed_gauss_blur_1_update_0_stage_165;
      bright_weights_normed_gauss_blur_1_update_0_stage_167 <= bright_weights_normed_gauss_blur_1_update_0_stage_166;
      bright_weights_normed_gauss_blur_1_update_0_stage_168 <= bright_weights_normed_gauss_blur_1_update_0_stage_167;
      bright_weights_normed_gauss_blur_1_update_0_stage_169 <= bright_weights_normed_gauss_blur_1_update_0_stage_168;
      bright_weights_normed_gauss_blur_1_update_0_stage_170 <= bright_weights_normed_gauss_blur_1_update_0_stage_169;
      bright_weights_normed_gauss_blur_1_update_0_stage_171 <= bright_weights_normed_gauss_blur_1_update_0_stage_170;
      bright_weights_normed_gauss_blur_1_update_0_stage_172 <= bright_weights_normed_gauss_blur_1_update_0_stage_171;
      bright_weights_normed_gauss_blur_1_update_0_stage_173 <= bright_weights_normed_gauss_blur_1_update_0_stage_172;
      bright_weights_normed_gauss_blur_1_update_0_stage_174 <= bright_weights_normed_gauss_blur_1_update_0_stage_173;
      bright_weights_normed_gauss_blur_1_update_0_stage_175 <= bright_weights_normed_gauss_blur_1_update_0_stage_174;
      bright_weights_normed_gauss_blur_1_update_0_stage_176 <= bright_weights_normed_gauss_blur_1_update_0_stage_175;
      bright_weights_normed_gauss_blur_1_update_0_stage_177 <= bright_weights_normed_gauss_blur_1_update_0_stage_176;
      bright_weights_normed_gauss_blur_1_update_0_stage_178 <= bright_weights_normed_gauss_blur_1_update_0_stage_177;
      bright_weights_normed_gauss_blur_1_update_0_stage_179 <= bright_weights_normed_gauss_blur_1_update_0_stage_178;
      bright_weights_normed_gauss_blur_1_update_0_stage_180 <= bright_weights_normed_gauss_blur_1_update_0_stage_179;
      bright_weights_normed_gauss_blur_1_update_0_stage_181 <= bright_weights_normed_gauss_blur_1_update_0_stage_180;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_82 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_83 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_82;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_84 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_83;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_85 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_84;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_86 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_85;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_87 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_86;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_88 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_87;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_89 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_88;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_90 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_89;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_91 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_90;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_92 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_91;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_93 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_92;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_94 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_93;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_95 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_94;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_96 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_95;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_97 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_96;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_98 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_97;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_99 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_98;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_100 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_99;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_101 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_100;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_102 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_101;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_103 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_102;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_104 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_103;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_105 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_104;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_106 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_105;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_107 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_106;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_108 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_107;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_109 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_108;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_110 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_109;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_111 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_110;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_112 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_111;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_113 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_112;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_114 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_113;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_115 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_114;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_116 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_115;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_117 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_116;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_118 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_117;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_119 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_118;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_120 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_119;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_121 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_120;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_122 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_121;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_123 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_122;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_124 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_123;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_125 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_124;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_126 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_125;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_127 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_126;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_128 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_127;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_129 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_128;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_130 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_129;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_131 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_130;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_132 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_131;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_133 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_132;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_134 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_133;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_135 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_134;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_136 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_135;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_137 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_136;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_138 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_137;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_139 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_138;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_140 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_139;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_141 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_140;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_142 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_141;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_143 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_142;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_144 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_143;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_145 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_144;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_146 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_145;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_147 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_146;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_148 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_147;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_149 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_148;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_150 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_149;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_151 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_150;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_152 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_151;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_153 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_152;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_154 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_153;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_155 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_154;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_156 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_155;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_157 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_156;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_158 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_157;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_159 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_158;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_160 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_159;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_161 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_160;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_162 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_161;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_163 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_162;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_164 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_163;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_165 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_164;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_166 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_165;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_167 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_166;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_168 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_167;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_169 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_168;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_170 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_169;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_171 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_170;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_172 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_171;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_173 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_172;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_174 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_173;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_175 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_174;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_176 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_175;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_177 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_176;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_178 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_177;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_179 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_178;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_180 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_179;
      bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_181 <= bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55_stage_180;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_88 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_89 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_88;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_90 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_89;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_91 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_90;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_92 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_91;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_93 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_92;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_94 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_93;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_95 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_94;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_96 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_95;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_97 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_96;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_98 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_97;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_99 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_98;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_100 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_99;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_101 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_100;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_102 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_101;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_103 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_102;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_104 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_103;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_105 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_104;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_106 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_105;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_107 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_106;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_108 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_107;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_109 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_108;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_110 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_109;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_111 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_110;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_112 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_111;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_113 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_112;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_114 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_113;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_115 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_114;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_116 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_115;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_117 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_116;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_118 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_117;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_119 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_118;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_120 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_119;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_121 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_120;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_122 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_121;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_123 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_122;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_124 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_123;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_125 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_124;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_126 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_125;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_127 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_126;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_128 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_127;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_129 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_128;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_130 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_129;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_131 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_130;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_132 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_131;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_133 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_132;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_134 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_133;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_135 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_134;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_136 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_135;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_137 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_136;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_138 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_137;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_139 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_138;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_140 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_139;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_141 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_140;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_142 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_141;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_143 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_142;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_144 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_143;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_145 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_144;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_146 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_145;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_147 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_146;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_148 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_147;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_149 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_148;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_150 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_149;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_151 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_150;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_152 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_151;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_153 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_152;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_154 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_153;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_155 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_154;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_156 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_155;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_157 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_156;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_158 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_157;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_159 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_158;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_160 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_159;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_161 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_160;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_162 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_161;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_163 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_162;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_164 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_163;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_165 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_164;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_166 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_165;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_167 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_166;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_168 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_167;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_169 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_168;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_170 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_169;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_171 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_170;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_172 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_171;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_173 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_172;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_174 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_173;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_175 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_174;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_176 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_175;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_177 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_176;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_178 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_177;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_179 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_178;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_180 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_179;
      bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_181 <= bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59_stage_180;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_84 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_85 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_84;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_86 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_85;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_87 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_86;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_88 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_87;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_89 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_88;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_90 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_89;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_91 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_90;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_92 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_91;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_93 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_92;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_94 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_93;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_95 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_94;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_96 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_95;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_97 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_96;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_98 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_97;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_99 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_98;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_100 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_99;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_101 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_100;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_102 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_101;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_103 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_102;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_104 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_103;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_105 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_104;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_106 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_105;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_107 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_106;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_108 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_107;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_109 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_108;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_110 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_109;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_111 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_110;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_112 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_111;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_113 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_112;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_114 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_113;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_115 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_114;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_116 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_115;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_117 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_116;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_118 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_117;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_119 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_118;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_120 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_119;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_121 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_120;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_122 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_121;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_123 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_122;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_124 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_123;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_125 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_124;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_126 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_125;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_127 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_126;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_128 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_127;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_129 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_128;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_130 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_129;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_131 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_130;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_132 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_131;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_133 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_132;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_134 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_133;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_135 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_134;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_136 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_135;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_137 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_136;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_138 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_137;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_139 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_138;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_140 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_139;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_141 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_140;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_142 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_141;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_143 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_142;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_144 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_143;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_145 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_144;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_146 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_145;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_147 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_146;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_148 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_147;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_149 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_148;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_150 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_149;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_151 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_150;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_152 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_151;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_153 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_152;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_154 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_153;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_155 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_154;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_156 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_155;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_157 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_156;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_158 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_157;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_159 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_158;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_160 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_159;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_161 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_160;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_162 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_161;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_163 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_162;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_164 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_163;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_165 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_164;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_166 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_165;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_167 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_166;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_168 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_167;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_169 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_168;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_170 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_169;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_171 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_170;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_172 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_171;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_173 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_172;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_174 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_173;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_175 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_174;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_176 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_175;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_177 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_176;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_178 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_177;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_179 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_178;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_180 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_179;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_181 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56_stage_180;
      bright_laplace_us_2_update_0_stage_89 <= bright_laplace_us_2_update_0;
      bright_laplace_us_2_update_0_stage_90 <= bright_laplace_us_2_update_0_stage_89;
      bright_laplace_us_2_update_0_stage_91 <= bright_laplace_us_2_update_0_stage_90;
      bright_laplace_us_2_update_0_stage_92 <= bright_laplace_us_2_update_0_stage_91;
      bright_laplace_us_2_update_0_stage_93 <= bright_laplace_us_2_update_0_stage_92;
      bright_laplace_us_2_update_0_stage_94 <= bright_laplace_us_2_update_0_stage_93;
      bright_laplace_us_2_update_0_stage_95 <= bright_laplace_us_2_update_0_stage_94;
      bright_laplace_us_2_update_0_stage_96 <= bright_laplace_us_2_update_0_stage_95;
      bright_laplace_us_2_update_0_stage_97 <= bright_laplace_us_2_update_0_stage_96;
      bright_laplace_us_2_update_0_stage_98 <= bright_laplace_us_2_update_0_stage_97;
      bright_laplace_us_2_update_0_stage_99 <= bright_laplace_us_2_update_0_stage_98;
      bright_laplace_us_2_update_0_stage_100 <= bright_laplace_us_2_update_0_stage_99;
      bright_laplace_us_2_update_0_stage_101 <= bright_laplace_us_2_update_0_stage_100;
      bright_laplace_us_2_update_0_stage_102 <= bright_laplace_us_2_update_0_stage_101;
      bright_laplace_us_2_update_0_stage_103 <= bright_laplace_us_2_update_0_stage_102;
      bright_laplace_us_2_update_0_stage_104 <= bright_laplace_us_2_update_0_stage_103;
      bright_laplace_us_2_update_0_stage_105 <= bright_laplace_us_2_update_0_stage_104;
      bright_laplace_us_2_update_0_stage_106 <= bright_laplace_us_2_update_0_stage_105;
      bright_laplace_us_2_update_0_stage_107 <= bright_laplace_us_2_update_0_stage_106;
      bright_laplace_us_2_update_0_stage_108 <= bright_laplace_us_2_update_0_stage_107;
      bright_laplace_us_2_update_0_stage_109 <= bright_laplace_us_2_update_0_stage_108;
      bright_laplace_us_2_update_0_stage_110 <= bright_laplace_us_2_update_0_stage_109;
      bright_laplace_us_2_update_0_stage_111 <= bright_laplace_us_2_update_0_stage_110;
      bright_laplace_us_2_update_0_stage_112 <= bright_laplace_us_2_update_0_stage_111;
      bright_laplace_us_2_update_0_stage_113 <= bright_laplace_us_2_update_0_stage_112;
      bright_laplace_us_2_update_0_stage_114 <= bright_laplace_us_2_update_0_stage_113;
      bright_laplace_us_2_update_0_stage_115 <= bright_laplace_us_2_update_0_stage_114;
      bright_laplace_us_2_update_0_stage_116 <= bright_laplace_us_2_update_0_stage_115;
      bright_laplace_us_2_update_0_stage_117 <= bright_laplace_us_2_update_0_stage_116;
      bright_laplace_us_2_update_0_stage_118 <= bright_laplace_us_2_update_0_stage_117;
      bright_laplace_us_2_update_0_stage_119 <= bright_laplace_us_2_update_0_stage_118;
      bright_laplace_us_2_update_0_stage_120 <= bright_laplace_us_2_update_0_stage_119;
      bright_laplace_us_2_update_0_stage_121 <= bright_laplace_us_2_update_0_stage_120;
      bright_laplace_us_2_update_0_stage_122 <= bright_laplace_us_2_update_0_stage_121;
      bright_laplace_us_2_update_0_stage_123 <= bright_laplace_us_2_update_0_stage_122;
      bright_laplace_us_2_update_0_stage_124 <= bright_laplace_us_2_update_0_stage_123;
      bright_laplace_us_2_update_0_stage_125 <= bright_laplace_us_2_update_0_stage_124;
      bright_laplace_us_2_update_0_stage_126 <= bright_laplace_us_2_update_0_stage_125;
      bright_laplace_us_2_update_0_stage_127 <= bright_laplace_us_2_update_0_stage_126;
      bright_laplace_us_2_update_0_stage_128 <= bright_laplace_us_2_update_0_stage_127;
      bright_laplace_us_2_update_0_stage_129 <= bright_laplace_us_2_update_0_stage_128;
      bright_laplace_us_2_update_0_stage_130 <= bright_laplace_us_2_update_0_stage_129;
      bright_laplace_us_2_update_0_stage_131 <= bright_laplace_us_2_update_0_stage_130;
      bright_laplace_us_2_update_0_stage_132 <= bright_laplace_us_2_update_0_stage_131;
      bright_laplace_us_2_update_0_stage_133 <= bright_laplace_us_2_update_0_stage_132;
      bright_laplace_us_2_update_0_stage_134 <= bright_laplace_us_2_update_0_stage_133;
      bright_laplace_us_2_update_0_stage_135 <= bright_laplace_us_2_update_0_stage_134;
      bright_laplace_us_2_update_0_stage_136 <= bright_laplace_us_2_update_0_stage_135;
      bright_laplace_us_2_update_0_stage_137 <= bright_laplace_us_2_update_0_stage_136;
      bright_laplace_us_2_update_0_stage_138 <= bright_laplace_us_2_update_0_stage_137;
      bright_laplace_us_2_update_0_stage_139 <= bright_laplace_us_2_update_0_stage_138;
      bright_laplace_us_2_update_0_stage_140 <= bright_laplace_us_2_update_0_stage_139;
      bright_laplace_us_2_update_0_stage_141 <= bright_laplace_us_2_update_0_stage_140;
      bright_laplace_us_2_update_0_stage_142 <= bright_laplace_us_2_update_0_stage_141;
      bright_laplace_us_2_update_0_stage_143 <= bright_laplace_us_2_update_0_stage_142;
      bright_laplace_us_2_update_0_stage_144 <= bright_laplace_us_2_update_0_stage_143;
      bright_laplace_us_2_update_0_stage_145 <= bright_laplace_us_2_update_0_stage_144;
      bright_laplace_us_2_update_0_stage_146 <= bright_laplace_us_2_update_0_stage_145;
      bright_laplace_us_2_update_0_stage_147 <= bright_laplace_us_2_update_0_stage_146;
      bright_laplace_us_2_update_0_stage_148 <= bright_laplace_us_2_update_0_stage_147;
      bright_laplace_us_2_update_0_stage_149 <= bright_laplace_us_2_update_0_stage_148;
      bright_laplace_us_2_update_0_stage_150 <= bright_laplace_us_2_update_0_stage_149;
      bright_laplace_us_2_update_0_stage_151 <= bright_laplace_us_2_update_0_stage_150;
      bright_laplace_us_2_update_0_stage_152 <= bright_laplace_us_2_update_0_stage_151;
      bright_laplace_us_2_update_0_stage_153 <= bright_laplace_us_2_update_0_stage_152;
      bright_laplace_us_2_update_0_stage_154 <= bright_laplace_us_2_update_0_stage_153;
      bright_laplace_us_2_update_0_stage_155 <= bright_laplace_us_2_update_0_stage_154;
      bright_laplace_us_2_update_0_stage_156 <= bright_laplace_us_2_update_0_stage_155;
      bright_laplace_us_2_update_0_stage_157 <= bright_laplace_us_2_update_0_stage_156;
      bright_laplace_us_2_update_0_stage_158 <= bright_laplace_us_2_update_0_stage_157;
      bright_laplace_us_2_update_0_stage_159 <= bright_laplace_us_2_update_0_stage_158;
      bright_laplace_us_2_update_0_stage_160 <= bright_laplace_us_2_update_0_stage_159;
      bright_laplace_us_2_update_0_stage_161 <= bright_laplace_us_2_update_0_stage_160;
      bright_laplace_us_2_update_0_stage_162 <= bright_laplace_us_2_update_0_stage_161;
      bright_laplace_us_2_update_0_stage_163 <= bright_laplace_us_2_update_0_stage_162;
      bright_laplace_us_2_update_0_stage_164 <= bright_laplace_us_2_update_0_stage_163;
      bright_laplace_us_2_update_0_stage_165 <= bright_laplace_us_2_update_0_stage_164;
      bright_laplace_us_2_update_0_stage_166 <= bright_laplace_us_2_update_0_stage_165;
      bright_laplace_us_2_update_0_stage_167 <= bright_laplace_us_2_update_0_stage_166;
      bright_laplace_us_2_update_0_stage_168 <= bright_laplace_us_2_update_0_stage_167;
      bright_laplace_us_2_update_0_stage_169 <= bright_laplace_us_2_update_0_stage_168;
      bright_laplace_us_2_update_0_stage_170 <= bright_laplace_us_2_update_0_stage_169;
      bright_laplace_us_2_update_0_stage_171 <= bright_laplace_us_2_update_0_stage_170;
      bright_laplace_us_2_update_0_stage_172 <= bright_laplace_us_2_update_0_stage_171;
      bright_laplace_us_2_update_0_stage_173 <= bright_laplace_us_2_update_0_stage_172;
      bright_laplace_us_2_update_0_stage_174 <= bright_laplace_us_2_update_0_stage_173;
      bright_laplace_us_2_update_0_stage_175 <= bright_laplace_us_2_update_0_stage_174;
      bright_laplace_us_2_update_0_stage_176 <= bright_laplace_us_2_update_0_stage_175;
      bright_laplace_us_2_update_0_stage_177 <= bright_laplace_us_2_update_0_stage_176;
      bright_laplace_us_2_update_0_stage_178 <= bright_laplace_us_2_update_0_stage_177;
      bright_laplace_us_2_update_0_stage_179 <= bright_laplace_us_2_update_0_stage_178;
      bright_laplace_us_2_update_0_stage_180 <= bright_laplace_us_2_update_0_stage_179;
      bright_laplace_us_2_update_0_stage_181 <= bright_laplace_us_2_update_0_stage_180;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_90 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_91 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_90;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_92 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_91;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_93 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_92;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_94 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_93;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_95 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_94;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_96 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_95;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_97 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_96;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_98 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_97;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_99 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_98;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_100 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_99;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_101 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_100;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_102 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_101;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_103 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_102;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_104 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_103;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_105 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_104;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_106 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_105;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_107 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_106;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_108 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_107;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_109 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_108;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_110 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_109;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_111 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_110;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_112 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_111;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_113 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_112;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_114 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_113;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_115 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_114;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_116 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_115;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_117 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_116;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_118 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_117;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_119 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_118;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_120 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_119;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_121 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_120;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_122 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_121;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_123 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_122;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_124 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_123;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_125 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_124;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_126 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_125;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_127 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_126;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_128 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_127;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_129 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_128;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_130 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_129;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_131 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_130;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_132 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_131;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_133 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_132;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_134 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_133;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_135 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_134;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_136 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_135;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_137 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_136;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_138 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_137;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_139 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_138;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_140 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_139;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_141 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_140;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_142 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_141;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_143 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_142;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_144 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_143;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_145 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_144;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_146 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_145;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_147 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_146;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_148 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_147;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_149 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_148;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_150 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_149;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_151 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_150;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_152 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_151;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_153 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_152;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_154 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_153;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_155 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_154;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_156 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_155;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_157 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_156;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_158 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_157;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_159 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_158;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_160 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_159;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_161 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_160;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_162 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_161;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_163 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_162;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_164 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_163;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_165 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_164;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_166 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_165;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_167 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_166;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_168 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_167;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_169 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_168;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_170 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_169;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_171 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_170;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_172 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_171;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_173 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_172;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_174 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_173;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_175 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_174;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_176 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_175;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_177 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_176;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_178 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_177;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_179 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_178;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_180 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_179;
      bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_181 <= bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60_stage_180;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_91 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_92 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_91;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_93 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_92;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_94 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_93;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_95 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_94;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_96 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_95;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_97 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_96;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_98 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_97;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_99 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_98;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_100 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_99;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_101 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_100;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_102 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_101;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_103 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_102;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_104 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_103;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_105 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_104;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_106 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_105;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_107 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_106;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_108 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_107;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_109 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_108;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_110 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_109;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_111 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_110;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_112 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_111;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_113 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_112;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_114 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_113;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_115 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_114;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_116 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_115;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_117 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_116;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_118 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_117;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_119 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_118;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_120 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_119;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_121 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_120;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_122 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_121;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_123 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_122;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_124 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_123;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_125 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_124;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_126 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_125;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_127 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_126;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_128 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_127;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_129 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_128;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_130 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_129;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_131 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_130;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_132 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_131;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_133 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_132;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_134 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_133;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_135 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_134;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_136 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_135;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_137 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_136;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_138 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_137;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_139 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_138;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_140 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_139;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_141 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_140;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_142 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_141;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_143 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_142;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_144 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_143;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_145 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_144;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_146 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_145;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_147 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_146;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_148 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_147;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_149 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_148;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_150 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_149;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_151 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_150;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_152 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_151;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_153 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_152;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_154 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_153;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_155 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_154;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_156 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_155;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_157 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_156;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_158 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_157;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_159 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_158;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_160 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_159;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_161 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_160;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_162 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_161;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_163 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_162;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_164 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_163;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_165 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_164;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_166 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_165;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_167 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_166;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_168 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_167;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_169 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_168;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_170 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_169;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_171 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_170;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_172 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_171;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_173 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_172;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_174 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_173;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_175 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_174;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_176 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_175;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_177 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_176;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_178 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_177;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_179 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_178;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_180 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_179;
      dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_181 <= dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61_stage_180;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_148 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_149 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_148;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_150 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_149;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_151 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_150;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_152 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_151;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_153 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_152;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_154 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_153;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_155 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_154;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_156 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_155;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_157 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_156;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_158 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_157;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_159 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_158;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_160 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_159;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_161 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_160;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_162 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_161;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_163 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_162;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_164 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_163;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_165 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_164;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_166 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_165;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_167 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_166;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_168 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_167;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_169 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_168;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_170 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_169;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_171 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_170;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_172 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_171;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_173 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_172;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_174 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_173;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_175 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_174;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_176 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_175;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_177 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_176;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_178 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_177;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_179 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_178;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_180 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_179;
      dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_181 <= dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102_stage_180;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_163 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_164 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_163;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_165 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_164;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_166 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_165;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_167 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_166;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_168 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_167;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_169 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_168;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_170 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_169;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_171 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_170;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_172 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_171;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_173 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_172;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_174 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_173;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_175 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_174;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_176 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_175;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_177 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_176;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_178 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_177;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_179 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_178;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_180 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_179;
      bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_181 <= bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114_stage_180;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_164 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_165 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_164;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_166 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_165;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_167 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_166;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_168 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_167;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_169 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_168;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_170 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_169;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_171 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_170;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_172 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_171;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_173 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_172;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_174 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_173;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_175 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_174;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_176 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_175;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_177 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_176;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_178 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_177;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_179 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_178;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_180 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_179;
      dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_181 <= dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115_stage_180;
      fused_level_3_update_0_stage_165 <= fused_level_3_update_0;
      fused_level_3_update_0_stage_166 <= fused_level_3_update_0_stage_165;
      fused_level_3_update_0_stage_167 <= fused_level_3_update_0_stage_166;
      fused_level_3_update_0_stage_168 <= fused_level_3_update_0_stage_167;
      fused_level_3_update_0_stage_169 <= fused_level_3_update_0_stage_168;
      fused_level_3_update_0_stage_170 <= fused_level_3_update_0_stage_169;
      fused_level_3_update_0_stage_171 <= fused_level_3_update_0_stage_170;
      fused_level_3_update_0_stage_172 <= fused_level_3_update_0_stage_171;
      fused_level_3_update_0_stage_173 <= fused_level_3_update_0_stage_172;
      fused_level_3_update_0_stage_174 <= fused_level_3_update_0_stage_173;
      fused_level_3_update_0_stage_175 <= fused_level_3_update_0_stage_174;
      fused_level_3_update_0_stage_176 <= fused_level_3_update_0_stage_175;
      fused_level_3_update_0_stage_177 <= fused_level_3_update_0_stage_176;
      fused_level_3_update_0_stage_178 <= fused_level_3_update_0_stage_177;
      fused_level_3_update_0_stage_179 <= fused_level_3_update_0_stage_178;
      fused_level_3_update_0_stage_180 <= fused_level_3_update_0_stage_179;
      fused_level_3_update_0_stage_181 <= fused_level_3_update_0_stage_180;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_166 <= fused_level_3_fused_level_3_update_0_write_write_116;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_167 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_166;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_168 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_167;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_169 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_168;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_170 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_169;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_171 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_170;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_172 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_171;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_173 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_172;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_174 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_173;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_175 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_174;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_176 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_175;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_177 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_176;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_178 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_177;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_179 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_178;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_180 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_179;
      fused_level_3_fused_level_3_update_0_write_write_116_stage_181 <= fused_level_3_fused_level_3_update_0_write_write_116_stage_180;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_167 <= fused_level_3_final_merged_2_update_0_read_read_117;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_168 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_167;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_169 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_168;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_170 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_169;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_171 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_170;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_172 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_171;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_173 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_172;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_174 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_173;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_175 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_174;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_176 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_175;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_177 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_176;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_178 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_177;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_179 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_178;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_180 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_179;
      fused_level_3_final_merged_2_update_0_read_read_117_stage_181 <= fused_level_3_final_merged_2_update_0_read_read_117_stage_180;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_168 <= fused_level_2_final_merged_2_update_0_read_read_118;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_169 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_168;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_170 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_169;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_171 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_170;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_172 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_171;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_173 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_172;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_174 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_173;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_175 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_174;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_176 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_175;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_177 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_176;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_178 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_177;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_179 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_178;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_180 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_179;
      fused_level_2_final_merged_2_update_0_read_read_118_stage_181 <= fused_level_2_final_merged_2_update_0_read_read_118_stage_180;
      final_merged_2_update_0_stage_169 <= final_merged_2_update_0;
      final_merged_2_update_0_stage_170 <= final_merged_2_update_0_stage_169;
      final_merged_2_update_0_stage_171 <= final_merged_2_update_0_stage_170;
      final_merged_2_update_0_stage_172 <= final_merged_2_update_0_stage_171;
      final_merged_2_update_0_stage_173 <= final_merged_2_update_0_stage_172;
      final_merged_2_update_0_stage_174 <= final_merged_2_update_0_stage_173;
      final_merged_2_update_0_stage_175 <= final_merged_2_update_0_stage_174;
      final_merged_2_update_0_stage_176 <= final_merged_2_update_0_stage_175;
      final_merged_2_update_0_stage_177 <= final_merged_2_update_0_stage_176;
      final_merged_2_update_0_stage_178 <= final_merged_2_update_0_stage_177;
      final_merged_2_update_0_stage_179 <= final_merged_2_update_0_stage_178;
      final_merged_2_update_0_stage_180 <= final_merged_2_update_0_stage_179;
      final_merged_2_update_0_stage_181 <= final_merged_2_update_0_stage_180;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_170 <= final_merged_2_final_merged_2_update_0_write_write_119;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_171 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_170;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_172 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_171;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_173 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_172;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_174 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_173;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_175 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_174;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_176 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_175;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_177 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_176;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_178 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_177;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_179 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_178;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_180 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_179;
      final_merged_2_final_merged_2_update_0_write_write_119_stage_181 <= final_merged_2_final_merged_2_update_0_write_write_119_stage_180;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_175 <= final_merged_1_final_merged_0_update_0_read_read_123;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_176 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_175;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_177 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_176;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_178 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_177;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_179 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_178;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_180 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_179;
      final_merged_1_final_merged_0_update_0_read_read_123_stage_181 <= final_merged_1_final_merged_0_update_0_read_read_123_stage_180;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_176 <= fused_level_0_final_merged_0_update_0_read_read_124;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_177 <= fused_level_0_final_merged_0_update_0_read_read_124_stage_176;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_178 <= fused_level_0_final_merged_0_update_0_read_read_124_stage_177;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_179 <= fused_level_0_final_merged_0_update_0_read_read_124_stage_178;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_180 <= fused_level_0_final_merged_0_update_0_read_read_124_stage_179;
      fused_level_0_final_merged_0_update_0_read_read_124_stage_181 <= fused_level_0_final_merged_0_update_0_read_read_124_stage_180;
      final_merged_0_update_0_stage_177 <= final_merged_0_update_0;
      final_merged_0_update_0_stage_178 <= final_merged_0_update_0_stage_177;
      final_merged_0_update_0_stage_179 <= final_merged_0_update_0_stage_178;
      final_merged_0_update_0_stage_180 <= final_merged_0_update_0_stage_179;
      final_merged_0_update_0_stage_181 <= final_merged_0_update_0_stage_180;
      final_merged_0_final_merged_0_update_0_write_write_125_stage_178 <= final_merged_0_final_merged_0_update_0_write_write_125;
      final_merged_0_final_merged_0_update_0_write_write_125_stage_179 <= final_merged_0_final_merged_0_update_0_write_write_125_stage_178;
      final_merged_0_final_merged_0_update_0_write_write_125_stage_180 <= final_merged_0_final_merged_0_update_0_write_write_125_stage_179;
      final_merged_0_final_merged_0_update_0_write_write_125_stage_181 <= final_merged_0_final_merged_0_update_0_write_write_125_stage_180;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_26 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_27 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_26;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_28 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_27;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_29 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_28;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_30 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_29;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_31 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_30;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_32 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_31;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_33 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_32;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_34 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_33;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_35 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_34;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_36 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_35;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_37 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_36;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_38 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_37;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_39 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_38;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_40 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_39;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_41 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_40;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_42 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_41;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_43 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_42;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_44 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_43;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_45 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_44;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_46 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_45;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_47 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_46;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_48 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_47;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_49 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_48;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_50 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_49;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_51 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_50;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_52 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_51;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_53 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_52;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_54 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_53;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_55 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_54;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_56 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_55;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_57 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_56;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_58 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_57;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_59 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_58;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_60 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_59;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_61 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_60;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_62 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_61;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_63 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_62;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_64 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_63;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_65 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_64;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_66 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_65;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_67 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_66;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_68 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_67;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_69 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_68;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_70 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_69;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_71 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_70;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_72 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_71;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_73 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_72;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_74 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_73;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_75 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_74;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_76 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_75;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_77 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_76;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_78 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_77;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_79 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_78;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_80 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_79;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_81 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_80;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_82 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_81;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_83 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_82;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_84 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_83;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_85 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_84;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_86 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_85;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_87 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_86;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_88 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_87;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_89 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_88;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_90 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_89;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_91 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_90;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_92 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_91;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_93 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_92;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_94 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_93;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_95 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_94;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_96 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_95;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_97 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_96;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_98 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_97;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_99 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_98;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_100 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_99;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_101 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_100;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_102 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_101;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_103 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_102;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_104 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_103;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_105 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_104;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_106 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_105;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_107 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_106;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_108 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_107;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_109 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_108;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_110 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_109;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_111 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_110;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_112 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_111;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_113 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_112;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_114 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_113;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_115 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_114;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_116 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_115;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_117 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_116;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_118 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_117;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_119 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_118;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_120 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_119;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_121 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_120;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_122 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_121;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_123 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_122;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_124 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_123;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_125 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_124;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_126 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_125;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_127 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_126;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_128 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_127;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_129 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_128;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_130 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_129;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_131 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_130;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_132 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_131;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_133 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_132;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_134 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_133;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_135 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_134;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_136 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_135;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_137 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_136;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_138 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_137;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_139 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_138;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_140 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_139;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_141 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_140;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_142 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_141;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_143 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_142;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_144 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_143;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_145 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_144;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_146 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_145;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_147 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_146;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_148 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_147;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_149 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_148;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_150 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_149;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_151 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_150;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_152 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_151;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_153 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_152;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_154 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_153;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_155 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_154;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_156 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_155;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_157 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_156;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_158 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_157;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_159 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_158;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_160 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_159;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_161 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_160;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_162 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_161;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_163 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_162;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_164 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_163;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_165 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_164;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_166 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_165;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_167 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_166;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_168 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_167;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_169 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_168;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_170 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_169;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_171 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_170;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_172 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_171;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_173 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_172;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_174 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_173;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_175 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_174;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_176 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_175;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_177 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_176;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_178 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_177;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_179 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_178;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_180 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_179;
      dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_181 <= dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16_stage_180;
      dark_laplace_us_0_update_0_stage_27 <= dark_laplace_us_0_update_0;
      dark_laplace_us_0_update_0_stage_28 <= dark_laplace_us_0_update_0_stage_27;
      dark_laplace_us_0_update_0_stage_29 <= dark_laplace_us_0_update_0_stage_28;
      dark_laplace_us_0_update_0_stage_30 <= dark_laplace_us_0_update_0_stage_29;
      dark_laplace_us_0_update_0_stage_31 <= dark_laplace_us_0_update_0_stage_30;
      dark_laplace_us_0_update_0_stage_32 <= dark_laplace_us_0_update_0_stage_31;
      dark_laplace_us_0_update_0_stage_33 <= dark_laplace_us_0_update_0_stage_32;
      dark_laplace_us_0_update_0_stage_34 <= dark_laplace_us_0_update_0_stage_33;
      dark_laplace_us_0_update_0_stage_35 <= dark_laplace_us_0_update_0_stage_34;
      dark_laplace_us_0_update_0_stage_36 <= dark_laplace_us_0_update_0_stage_35;
      dark_laplace_us_0_update_0_stage_37 <= dark_laplace_us_0_update_0_stage_36;
      dark_laplace_us_0_update_0_stage_38 <= dark_laplace_us_0_update_0_stage_37;
      dark_laplace_us_0_update_0_stage_39 <= dark_laplace_us_0_update_0_stage_38;
      dark_laplace_us_0_update_0_stage_40 <= dark_laplace_us_0_update_0_stage_39;
      dark_laplace_us_0_update_0_stage_41 <= dark_laplace_us_0_update_0_stage_40;
      dark_laplace_us_0_update_0_stage_42 <= dark_laplace_us_0_update_0_stage_41;
      dark_laplace_us_0_update_0_stage_43 <= dark_laplace_us_0_update_0_stage_42;
      dark_laplace_us_0_update_0_stage_44 <= dark_laplace_us_0_update_0_stage_43;
      dark_laplace_us_0_update_0_stage_45 <= dark_laplace_us_0_update_0_stage_44;
      dark_laplace_us_0_update_0_stage_46 <= dark_laplace_us_0_update_0_stage_45;
      dark_laplace_us_0_update_0_stage_47 <= dark_laplace_us_0_update_0_stage_46;
      dark_laplace_us_0_update_0_stage_48 <= dark_laplace_us_0_update_0_stage_47;
      dark_laplace_us_0_update_0_stage_49 <= dark_laplace_us_0_update_0_stage_48;
      dark_laplace_us_0_update_0_stage_50 <= dark_laplace_us_0_update_0_stage_49;
      dark_laplace_us_0_update_0_stage_51 <= dark_laplace_us_0_update_0_stage_50;
      dark_laplace_us_0_update_0_stage_52 <= dark_laplace_us_0_update_0_stage_51;
      dark_laplace_us_0_update_0_stage_53 <= dark_laplace_us_0_update_0_stage_52;
      dark_laplace_us_0_update_0_stage_54 <= dark_laplace_us_0_update_0_stage_53;
      dark_laplace_us_0_update_0_stage_55 <= dark_laplace_us_0_update_0_stage_54;
      dark_laplace_us_0_update_0_stage_56 <= dark_laplace_us_0_update_0_stage_55;
      dark_laplace_us_0_update_0_stage_57 <= dark_laplace_us_0_update_0_stage_56;
      dark_laplace_us_0_update_0_stage_58 <= dark_laplace_us_0_update_0_stage_57;
      dark_laplace_us_0_update_0_stage_59 <= dark_laplace_us_0_update_0_stage_58;
      dark_laplace_us_0_update_0_stage_60 <= dark_laplace_us_0_update_0_stage_59;
      dark_laplace_us_0_update_0_stage_61 <= dark_laplace_us_0_update_0_stage_60;
      dark_laplace_us_0_update_0_stage_62 <= dark_laplace_us_0_update_0_stage_61;
      dark_laplace_us_0_update_0_stage_63 <= dark_laplace_us_0_update_0_stage_62;
      dark_laplace_us_0_update_0_stage_64 <= dark_laplace_us_0_update_0_stage_63;
      dark_laplace_us_0_update_0_stage_65 <= dark_laplace_us_0_update_0_stage_64;
      dark_laplace_us_0_update_0_stage_66 <= dark_laplace_us_0_update_0_stage_65;
      dark_laplace_us_0_update_0_stage_67 <= dark_laplace_us_0_update_0_stage_66;
      dark_laplace_us_0_update_0_stage_68 <= dark_laplace_us_0_update_0_stage_67;
      dark_laplace_us_0_update_0_stage_69 <= dark_laplace_us_0_update_0_stage_68;
      dark_laplace_us_0_update_0_stage_70 <= dark_laplace_us_0_update_0_stage_69;
      dark_laplace_us_0_update_0_stage_71 <= dark_laplace_us_0_update_0_stage_70;
      dark_laplace_us_0_update_0_stage_72 <= dark_laplace_us_0_update_0_stage_71;
      dark_laplace_us_0_update_0_stage_73 <= dark_laplace_us_0_update_0_stage_72;
      dark_laplace_us_0_update_0_stage_74 <= dark_laplace_us_0_update_0_stage_73;
      dark_laplace_us_0_update_0_stage_75 <= dark_laplace_us_0_update_0_stage_74;
      dark_laplace_us_0_update_0_stage_76 <= dark_laplace_us_0_update_0_stage_75;
      dark_laplace_us_0_update_0_stage_77 <= dark_laplace_us_0_update_0_stage_76;
      dark_laplace_us_0_update_0_stage_78 <= dark_laplace_us_0_update_0_stage_77;
      dark_laplace_us_0_update_0_stage_79 <= dark_laplace_us_0_update_0_stage_78;
      dark_laplace_us_0_update_0_stage_80 <= dark_laplace_us_0_update_0_stage_79;
      dark_laplace_us_0_update_0_stage_81 <= dark_laplace_us_0_update_0_stage_80;
      dark_laplace_us_0_update_0_stage_82 <= dark_laplace_us_0_update_0_stage_81;
      dark_laplace_us_0_update_0_stage_83 <= dark_laplace_us_0_update_0_stage_82;
      dark_laplace_us_0_update_0_stage_84 <= dark_laplace_us_0_update_0_stage_83;
      dark_laplace_us_0_update_0_stage_85 <= dark_laplace_us_0_update_0_stage_84;
      dark_laplace_us_0_update_0_stage_86 <= dark_laplace_us_0_update_0_stage_85;
      dark_laplace_us_0_update_0_stage_87 <= dark_laplace_us_0_update_0_stage_86;
      dark_laplace_us_0_update_0_stage_88 <= dark_laplace_us_0_update_0_stage_87;
      dark_laplace_us_0_update_0_stage_89 <= dark_laplace_us_0_update_0_stage_88;
      dark_laplace_us_0_update_0_stage_90 <= dark_laplace_us_0_update_0_stage_89;
      dark_laplace_us_0_update_0_stage_91 <= dark_laplace_us_0_update_0_stage_90;
      dark_laplace_us_0_update_0_stage_92 <= dark_laplace_us_0_update_0_stage_91;
      dark_laplace_us_0_update_0_stage_93 <= dark_laplace_us_0_update_0_stage_92;
      dark_laplace_us_0_update_0_stage_94 <= dark_laplace_us_0_update_0_stage_93;
      dark_laplace_us_0_update_0_stage_95 <= dark_laplace_us_0_update_0_stage_94;
      dark_laplace_us_0_update_0_stage_96 <= dark_laplace_us_0_update_0_stage_95;
      dark_laplace_us_0_update_0_stage_97 <= dark_laplace_us_0_update_0_stage_96;
      dark_laplace_us_0_update_0_stage_98 <= dark_laplace_us_0_update_0_stage_97;
      dark_laplace_us_0_update_0_stage_99 <= dark_laplace_us_0_update_0_stage_98;
      dark_laplace_us_0_update_0_stage_100 <= dark_laplace_us_0_update_0_stage_99;
      dark_laplace_us_0_update_0_stage_101 <= dark_laplace_us_0_update_0_stage_100;
      dark_laplace_us_0_update_0_stage_102 <= dark_laplace_us_0_update_0_stage_101;
      dark_laplace_us_0_update_0_stage_103 <= dark_laplace_us_0_update_0_stage_102;
      dark_laplace_us_0_update_0_stage_104 <= dark_laplace_us_0_update_0_stage_103;
      dark_laplace_us_0_update_0_stage_105 <= dark_laplace_us_0_update_0_stage_104;
      dark_laplace_us_0_update_0_stage_106 <= dark_laplace_us_0_update_0_stage_105;
      dark_laplace_us_0_update_0_stage_107 <= dark_laplace_us_0_update_0_stage_106;
      dark_laplace_us_0_update_0_stage_108 <= dark_laplace_us_0_update_0_stage_107;
      dark_laplace_us_0_update_0_stage_109 <= dark_laplace_us_0_update_0_stage_108;
      dark_laplace_us_0_update_0_stage_110 <= dark_laplace_us_0_update_0_stage_109;
      dark_laplace_us_0_update_0_stage_111 <= dark_laplace_us_0_update_0_stage_110;
      dark_laplace_us_0_update_0_stage_112 <= dark_laplace_us_0_update_0_stage_111;
      dark_laplace_us_0_update_0_stage_113 <= dark_laplace_us_0_update_0_stage_112;
      dark_laplace_us_0_update_0_stage_114 <= dark_laplace_us_0_update_0_stage_113;
      dark_laplace_us_0_update_0_stage_115 <= dark_laplace_us_0_update_0_stage_114;
      dark_laplace_us_0_update_0_stage_116 <= dark_laplace_us_0_update_0_stage_115;
      dark_laplace_us_0_update_0_stage_117 <= dark_laplace_us_0_update_0_stage_116;
      dark_laplace_us_0_update_0_stage_118 <= dark_laplace_us_0_update_0_stage_117;
      dark_laplace_us_0_update_0_stage_119 <= dark_laplace_us_0_update_0_stage_118;
      dark_laplace_us_0_update_0_stage_120 <= dark_laplace_us_0_update_0_stage_119;
      dark_laplace_us_0_update_0_stage_121 <= dark_laplace_us_0_update_0_stage_120;
      dark_laplace_us_0_update_0_stage_122 <= dark_laplace_us_0_update_0_stage_121;
      dark_laplace_us_0_update_0_stage_123 <= dark_laplace_us_0_update_0_stage_122;
      dark_laplace_us_0_update_0_stage_124 <= dark_laplace_us_0_update_0_stage_123;
      dark_laplace_us_0_update_0_stage_125 <= dark_laplace_us_0_update_0_stage_124;
      dark_laplace_us_0_update_0_stage_126 <= dark_laplace_us_0_update_0_stage_125;
      dark_laplace_us_0_update_0_stage_127 <= dark_laplace_us_0_update_0_stage_126;
      dark_laplace_us_0_update_0_stage_128 <= dark_laplace_us_0_update_0_stage_127;
      dark_laplace_us_0_update_0_stage_129 <= dark_laplace_us_0_update_0_stage_128;
      dark_laplace_us_0_update_0_stage_130 <= dark_laplace_us_0_update_0_stage_129;
      dark_laplace_us_0_update_0_stage_131 <= dark_laplace_us_0_update_0_stage_130;
      dark_laplace_us_0_update_0_stage_132 <= dark_laplace_us_0_update_0_stage_131;
      dark_laplace_us_0_update_0_stage_133 <= dark_laplace_us_0_update_0_stage_132;
      dark_laplace_us_0_update_0_stage_134 <= dark_laplace_us_0_update_0_stage_133;
      dark_laplace_us_0_update_0_stage_135 <= dark_laplace_us_0_update_0_stage_134;
      dark_laplace_us_0_update_0_stage_136 <= dark_laplace_us_0_update_0_stage_135;
      dark_laplace_us_0_update_0_stage_137 <= dark_laplace_us_0_update_0_stage_136;
      dark_laplace_us_0_update_0_stage_138 <= dark_laplace_us_0_update_0_stage_137;
      dark_laplace_us_0_update_0_stage_139 <= dark_laplace_us_0_update_0_stage_138;
      dark_laplace_us_0_update_0_stage_140 <= dark_laplace_us_0_update_0_stage_139;
      dark_laplace_us_0_update_0_stage_141 <= dark_laplace_us_0_update_0_stage_140;
      dark_laplace_us_0_update_0_stage_142 <= dark_laplace_us_0_update_0_stage_141;
      dark_laplace_us_0_update_0_stage_143 <= dark_laplace_us_0_update_0_stage_142;
      dark_laplace_us_0_update_0_stage_144 <= dark_laplace_us_0_update_0_stage_143;
      dark_laplace_us_0_update_0_stage_145 <= dark_laplace_us_0_update_0_stage_144;
      dark_laplace_us_0_update_0_stage_146 <= dark_laplace_us_0_update_0_stage_145;
      dark_laplace_us_0_update_0_stage_147 <= dark_laplace_us_0_update_0_stage_146;
      dark_laplace_us_0_update_0_stage_148 <= dark_laplace_us_0_update_0_stage_147;
      dark_laplace_us_0_update_0_stage_149 <= dark_laplace_us_0_update_0_stage_148;
      dark_laplace_us_0_update_0_stage_150 <= dark_laplace_us_0_update_0_stage_149;
      dark_laplace_us_0_update_0_stage_151 <= dark_laplace_us_0_update_0_stage_150;
      dark_laplace_us_0_update_0_stage_152 <= dark_laplace_us_0_update_0_stage_151;
      dark_laplace_us_0_update_0_stage_153 <= dark_laplace_us_0_update_0_stage_152;
      dark_laplace_us_0_update_0_stage_154 <= dark_laplace_us_0_update_0_stage_153;
      dark_laplace_us_0_update_0_stage_155 <= dark_laplace_us_0_update_0_stage_154;
      dark_laplace_us_0_update_0_stage_156 <= dark_laplace_us_0_update_0_stage_155;
      dark_laplace_us_0_update_0_stage_157 <= dark_laplace_us_0_update_0_stage_156;
      dark_laplace_us_0_update_0_stage_158 <= dark_laplace_us_0_update_0_stage_157;
      dark_laplace_us_0_update_0_stage_159 <= dark_laplace_us_0_update_0_stage_158;
      dark_laplace_us_0_update_0_stage_160 <= dark_laplace_us_0_update_0_stage_159;
      dark_laplace_us_0_update_0_stage_161 <= dark_laplace_us_0_update_0_stage_160;
      dark_laplace_us_0_update_0_stage_162 <= dark_laplace_us_0_update_0_stage_161;
      dark_laplace_us_0_update_0_stage_163 <= dark_laplace_us_0_update_0_stage_162;
      dark_laplace_us_0_update_0_stage_164 <= dark_laplace_us_0_update_0_stage_163;
      dark_laplace_us_0_update_0_stage_165 <= dark_laplace_us_0_update_0_stage_164;
      dark_laplace_us_0_update_0_stage_166 <= dark_laplace_us_0_update_0_stage_165;
      dark_laplace_us_0_update_0_stage_167 <= dark_laplace_us_0_update_0_stage_166;
      dark_laplace_us_0_update_0_stage_168 <= dark_laplace_us_0_update_0_stage_167;
      dark_laplace_us_0_update_0_stage_169 <= dark_laplace_us_0_update_0_stage_168;
      dark_laplace_us_0_update_0_stage_170 <= dark_laplace_us_0_update_0_stage_169;
      dark_laplace_us_0_update_0_stage_171 <= dark_laplace_us_0_update_0_stage_170;
      dark_laplace_us_0_update_0_stage_172 <= dark_laplace_us_0_update_0_stage_171;
      dark_laplace_us_0_update_0_stage_173 <= dark_laplace_us_0_update_0_stage_172;
      dark_laplace_us_0_update_0_stage_174 <= dark_laplace_us_0_update_0_stage_173;
      dark_laplace_us_0_update_0_stage_175 <= dark_laplace_us_0_update_0_stage_174;
      dark_laplace_us_0_update_0_stage_176 <= dark_laplace_us_0_update_0_stage_175;
      dark_laplace_us_0_update_0_stage_177 <= dark_laplace_us_0_update_0_stage_176;
      dark_laplace_us_0_update_0_stage_178 <= dark_laplace_us_0_update_0_stage_177;
      dark_laplace_us_0_update_0_stage_179 <= dark_laplace_us_0_update_0_stage_178;
      dark_laplace_us_0_update_0_stage_180 <= dark_laplace_us_0_update_0_stage_179;
      dark_laplace_us_0_update_0_stage_181 <= dark_laplace_us_0_update_0_stage_180;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_28 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_29 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_28;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_30 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_29;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_31 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_30;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_32 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_31;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_33 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_32;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_34 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_33;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_35 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_34;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_36 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_35;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_37 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_36;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_38 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_37;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_39 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_38;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_40 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_39;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_41 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_40;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_42 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_41;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_43 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_42;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_44 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_43;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_45 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_44;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_46 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_45;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_47 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_46;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_48 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_47;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_49 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_48;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_50 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_49;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_51 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_50;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_52 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_51;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_53 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_52;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_54 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_53;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_55 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_54;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_56 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_55;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_57 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_56;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_58 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_57;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_59 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_58;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_60 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_59;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_61 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_60;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_62 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_61;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_63 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_62;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_64 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_63;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_65 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_64;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_66 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_65;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_67 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_66;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_68 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_67;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_69 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_68;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_70 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_69;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_71 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_70;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_72 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_71;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_73 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_72;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_74 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_73;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_75 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_74;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_76 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_75;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_77 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_76;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_78 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_77;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_79 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_78;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_80 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_79;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_81 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_80;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_82 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_81;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_83 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_82;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_84 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_83;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_85 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_84;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_86 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_85;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_87 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_86;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_88 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_87;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_89 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_88;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_90 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_89;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_91 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_90;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_92 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_91;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_93 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_92;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_94 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_93;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_95 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_94;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_96 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_95;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_97 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_96;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_98 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_97;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_99 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_98;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_100 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_99;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_101 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_100;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_102 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_101;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_103 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_102;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_104 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_103;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_105 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_104;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_106 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_105;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_107 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_106;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_108 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_107;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_109 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_108;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_110 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_109;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_111 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_110;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_112 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_111;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_113 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_112;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_114 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_113;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_115 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_114;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_116 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_115;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_117 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_116;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_118 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_117;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_119 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_118;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_120 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_119;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_121 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_120;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_122 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_121;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_123 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_122;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_124 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_123;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_125 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_124;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_126 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_125;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_127 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_126;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_128 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_127;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_129 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_128;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_130 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_129;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_131 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_130;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_132 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_131;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_133 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_132;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_134 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_133;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_135 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_134;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_136 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_135;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_137 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_136;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_138 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_137;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_139 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_138;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_140 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_139;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_141 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_140;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_142 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_141;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_143 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_142;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_144 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_143;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_145 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_144;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_146 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_145;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_147 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_146;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_148 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_147;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_149 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_148;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_150 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_149;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_151 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_150;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_152 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_151;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_153 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_152;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_154 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_153;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_155 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_154;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_156 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_155;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_157 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_156;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_158 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_157;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_159 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_158;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_160 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_159;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_161 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_160;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_162 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_161;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_163 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_162;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_164 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_163;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_165 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_164;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_166 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_165;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_167 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_166;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_168 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_167;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_169 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_168;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_170 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_169;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_171 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_170;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_172 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_171;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_173 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_172;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_174 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_173;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_175 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_174;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_176 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_175;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_177 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_176;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_178 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_177;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_179 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_178;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_180 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_179;
      dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_181 <= dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17_stage_180;
      dark_weights_weight_sums_update_0_read_read_22_stage_35 <= dark_weights_weight_sums_update_0_read_read_22;
      dark_weights_weight_sums_update_0_read_read_22_stage_36 <= dark_weights_weight_sums_update_0_read_read_22_stage_35;
      dark_weights_weight_sums_update_0_read_read_22_stage_37 <= dark_weights_weight_sums_update_0_read_read_22_stage_36;
      dark_weights_weight_sums_update_0_read_read_22_stage_38 <= dark_weights_weight_sums_update_0_read_read_22_stage_37;
      dark_weights_weight_sums_update_0_read_read_22_stage_39 <= dark_weights_weight_sums_update_0_read_read_22_stage_38;
      dark_weights_weight_sums_update_0_read_read_22_stage_40 <= dark_weights_weight_sums_update_0_read_read_22_stage_39;
      dark_weights_weight_sums_update_0_read_read_22_stage_41 <= dark_weights_weight_sums_update_0_read_read_22_stage_40;
      dark_weights_weight_sums_update_0_read_read_22_stage_42 <= dark_weights_weight_sums_update_0_read_read_22_stage_41;
      dark_weights_weight_sums_update_0_read_read_22_stage_43 <= dark_weights_weight_sums_update_0_read_read_22_stage_42;
      dark_weights_weight_sums_update_0_read_read_22_stage_44 <= dark_weights_weight_sums_update_0_read_read_22_stage_43;
      dark_weights_weight_sums_update_0_read_read_22_stage_45 <= dark_weights_weight_sums_update_0_read_read_22_stage_44;
      dark_weights_weight_sums_update_0_read_read_22_stage_46 <= dark_weights_weight_sums_update_0_read_read_22_stage_45;
      dark_weights_weight_sums_update_0_read_read_22_stage_47 <= dark_weights_weight_sums_update_0_read_read_22_stage_46;
      dark_weights_weight_sums_update_0_read_read_22_stage_48 <= dark_weights_weight_sums_update_0_read_read_22_stage_47;
      dark_weights_weight_sums_update_0_read_read_22_stage_49 <= dark_weights_weight_sums_update_0_read_read_22_stage_48;
      dark_weights_weight_sums_update_0_read_read_22_stage_50 <= dark_weights_weight_sums_update_0_read_read_22_stage_49;
      dark_weights_weight_sums_update_0_read_read_22_stage_51 <= dark_weights_weight_sums_update_0_read_read_22_stage_50;
      dark_weights_weight_sums_update_0_read_read_22_stage_52 <= dark_weights_weight_sums_update_0_read_read_22_stage_51;
      dark_weights_weight_sums_update_0_read_read_22_stage_53 <= dark_weights_weight_sums_update_0_read_read_22_stage_52;
      dark_weights_weight_sums_update_0_read_read_22_stage_54 <= dark_weights_weight_sums_update_0_read_read_22_stage_53;
      dark_weights_weight_sums_update_0_read_read_22_stage_55 <= dark_weights_weight_sums_update_0_read_read_22_stage_54;
      dark_weights_weight_sums_update_0_read_read_22_stage_56 <= dark_weights_weight_sums_update_0_read_read_22_stage_55;
      dark_weights_weight_sums_update_0_read_read_22_stage_57 <= dark_weights_weight_sums_update_0_read_read_22_stage_56;
      dark_weights_weight_sums_update_0_read_read_22_stage_58 <= dark_weights_weight_sums_update_0_read_read_22_stage_57;
      dark_weights_weight_sums_update_0_read_read_22_stage_59 <= dark_weights_weight_sums_update_0_read_read_22_stage_58;
      dark_weights_weight_sums_update_0_read_read_22_stage_60 <= dark_weights_weight_sums_update_0_read_read_22_stage_59;
      dark_weights_weight_sums_update_0_read_read_22_stage_61 <= dark_weights_weight_sums_update_0_read_read_22_stage_60;
      dark_weights_weight_sums_update_0_read_read_22_stage_62 <= dark_weights_weight_sums_update_0_read_read_22_stage_61;
      dark_weights_weight_sums_update_0_read_read_22_stage_63 <= dark_weights_weight_sums_update_0_read_read_22_stage_62;
      dark_weights_weight_sums_update_0_read_read_22_stage_64 <= dark_weights_weight_sums_update_0_read_read_22_stage_63;
      dark_weights_weight_sums_update_0_read_read_22_stage_65 <= dark_weights_weight_sums_update_0_read_read_22_stage_64;
      dark_weights_weight_sums_update_0_read_read_22_stage_66 <= dark_weights_weight_sums_update_0_read_read_22_stage_65;
      dark_weights_weight_sums_update_0_read_read_22_stage_67 <= dark_weights_weight_sums_update_0_read_read_22_stage_66;
      dark_weights_weight_sums_update_0_read_read_22_stage_68 <= dark_weights_weight_sums_update_0_read_read_22_stage_67;
      dark_weights_weight_sums_update_0_read_read_22_stage_69 <= dark_weights_weight_sums_update_0_read_read_22_stage_68;
      dark_weights_weight_sums_update_0_read_read_22_stage_70 <= dark_weights_weight_sums_update_0_read_read_22_stage_69;
      dark_weights_weight_sums_update_0_read_read_22_stage_71 <= dark_weights_weight_sums_update_0_read_read_22_stage_70;
      dark_weights_weight_sums_update_0_read_read_22_stage_72 <= dark_weights_weight_sums_update_0_read_read_22_stage_71;
      dark_weights_weight_sums_update_0_read_read_22_stage_73 <= dark_weights_weight_sums_update_0_read_read_22_stage_72;
      dark_weights_weight_sums_update_0_read_read_22_stage_74 <= dark_weights_weight_sums_update_0_read_read_22_stage_73;
      dark_weights_weight_sums_update_0_read_read_22_stage_75 <= dark_weights_weight_sums_update_0_read_read_22_stage_74;
      dark_weights_weight_sums_update_0_read_read_22_stage_76 <= dark_weights_weight_sums_update_0_read_read_22_stage_75;
      dark_weights_weight_sums_update_0_read_read_22_stage_77 <= dark_weights_weight_sums_update_0_read_read_22_stage_76;
      dark_weights_weight_sums_update_0_read_read_22_stage_78 <= dark_weights_weight_sums_update_0_read_read_22_stage_77;
      dark_weights_weight_sums_update_0_read_read_22_stage_79 <= dark_weights_weight_sums_update_0_read_read_22_stage_78;
      dark_weights_weight_sums_update_0_read_read_22_stage_80 <= dark_weights_weight_sums_update_0_read_read_22_stage_79;
      dark_weights_weight_sums_update_0_read_read_22_stage_81 <= dark_weights_weight_sums_update_0_read_read_22_stage_80;
      dark_weights_weight_sums_update_0_read_read_22_stage_82 <= dark_weights_weight_sums_update_0_read_read_22_stage_81;
      dark_weights_weight_sums_update_0_read_read_22_stage_83 <= dark_weights_weight_sums_update_0_read_read_22_stage_82;
      dark_weights_weight_sums_update_0_read_read_22_stage_84 <= dark_weights_weight_sums_update_0_read_read_22_stage_83;
      dark_weights_weight_sums_update_0_read_read_22_stage_85 <= dark_weights_weight_sums_update_0_read_read_22_stage_84;
      dark_weights_weight_sums_update_0_read_read_22_stage_86 <= dark_weights_weight_sums_update_0_read_read_22_stage_85;
      dark_weights_weight_sums_update_0_read_read_22_stage_87 <= dark_weights_weight_sums_update_0_read_read_22_stage_86;
      dark_weights_weight_sums_update_0_read_read_22_stage_88 <= dark_weights_weight_sums_update_0_read_read_22_stage_87;
      dark_weights_weight_sums_update_0_read_read_22_stage_89 <= dark_weights_weight_sums_update_0_read_read_22_stage_88;
      dark_weights_weight_sums_update_0_read_read_22_stage_90 <= dark_weights_weight_sums_update_0_read_read_22_stage_89;
      dark_weights_weight_sums_update_0_read_read_22_stage_91 <= dark_weights_weight_sums_update_0_read_read_22_stage_90;
      dark_weights_weight_sums_update_0_read_read_22_stage_92 <= dark_weights_weight_sums_update_0_read_read_22_stage_91;
      dark_weights_weight_sums_update_0_read_read_22_stage_93 <= dark_weights_weight_sums_update_0_read_read_22_stage_92;
      dark_weights_weight_sums_update_0_read_read_22_stage_94 <= dark_weights_weight_sums_update_0_read_read_22_stage_93;
      dark_weights_weight_sums_update_0_read_read_22_stage_95 <= dark_weights_weight_sums_update_0_read_read_22_stage_94;
      dark_weights_weight_sums_update_0_read_read_22_stage_96 <= dark_weights_weight_sums_update_0_read_read_22_stage_95;
      dark_weights_weight_sums_update_0_read_read_22_stage_97 <= dark_weights_weight_sums_update_0_read_read_22_stage_96;
      dark_weights_weight_sums_update_0_read_read_22_stage_98 <= dark_weights_weight_sums_update_0_read_read_22_stage_97;
      dark_weights_weight_sums_update_0_read_read_22_stage_99 <= dark_weights_weight_sums_update_0_read_read_22_stage_98;
      dark_weights_weight_sums_update_0_read_read_22_stage_100 <= dark_weights_weight_sums_update_0_read_read_22_stage_99;
      dark_weights_weight_sums_update_0_read_read_22_stage_101 <= dark_weights_weight_sums_update_0_read_read_22_stage_100;
      dark_weights_weight_sums_update_0_read_read_22_stage_102 <= dark_weights_weight_sums_update_0_read_read_22_stage_101;
      dark_weights_weight_sums_update_0_read_read_22_stage_103 <= dark_weights_weight_sums_update_0_read_read_22_stage_102;
      dark_weights_weight_sums_update_0_read_read_22_stage_104 <= dark_weights_weight_sums_update_0_read_read_22_stage_103;
      dark_weights_weight_sums_update_0_read_read_22_stage_105 <= dark_weights_weight_sums_update_0_read_read_22_stage_104;
      dark_weights_weight_sums_update_0_read_read_22_stage_106 <= dark_weights_weight_sums_update_0_read_read_22_stage_105;
      dark_weights_weight_sums_update_0_read_read_22_stage_107 <= dark_weights_weight_sums_update_0_read_read_22_stage_106;
      dark_weights_weight_sums_update_0_read_read_22_stage_108 <= dark_weights_weight_sums_update_0_read_read_22_stage_107;
      dark_weights_weight_sums_update_0_read_read_22_stage_109 <= dark_weights_weight_sums_update_0_read_read_22_stage_108;
      dark_weights_weight_sums_update_0_read_read_22_stage_110 <= dark_weights_weight_sums_update_0_read_read_22_stage_109;
      dark_weights_weight_sums_update_0_read_read_22_stage_111 <= dark_weights_weight_sums_update_0_read_read_22_stage_110;
      dark_weights_weight_sums_update_0_read_read_22_stage_112 <= dark_weights_weight_sums_update_0_read_read_22_stage_111;
      dark_weights_weight_sums_update_0_read_read_22_stage_113 <= dark_weights_weight_sums_update_0_read_read_22_stage_112;
      dark_weights_weight_sums_update_0_read_read_22_stage_114 <= dark_weights_weight_sums_update_0_read_read_22_stage_113;
      dark_weights_weight_sums_update_0_read_read_22_stage_115 <= dark_weights_weight_sums_update_0_read_read_22_stage_114;
      dark_weights_weight_sums_update_0_read_read_22_stage_116 <= dark_weights_weight_sums_update_0_read_read_22_stage_115;
      dark_weights_weight_sums_update_0_read_read_22_stage_117 <= dark_weights_weight_sums_update_0_read_read_22_stage_116;
      dark_weights_weight_sums_update_0_read_read_22_stage_118 <= dark_weights_weight_sums_update_0_read_read_22_stage_117;
      dark_weights_weight_sums_update_0_read_read_22_stage_119 <= dark_weights_weight_sums_update_0_read_read_22_stage_118;
      dark_weights_weight_sums_update_0_read_read_22_stage_120 <= dark_weights_weight_sums_update_0_read_read_22_stage_119;
      dark_weights_weight_sums_update_0_read_read_22_stage_121 <= dark_weights_weight_sums_update_0_read_read_22_stage_120;
      dark_weights_weight_sums_update_0_read_read_22_stage_122 <= dark_weights_weight_sums_update_0_read_read_22_stage_121;
      dark_weights_weight_sums_update_0_read_read_22_stage_123 <= dark_weights_weight_sums_update_0_read_read_22_stage_122;
      dark_weights_weight_sums_update_0_read_read_22_stage_124 <= dark_weights_weight_sums_update_0_read_read_22_stage_123;
      dark_weights_weight_sums_update_0_read_read_22_stage_125 <= dark_weights_weight_sums_update_0_read_read_22_stage_124;
      dark_weights_weight_sums_update_0_read_read_22_stage_126 <= dark_weights_weight_sums_update_0_read_read_22_stage_125;
      dark_weights_weight_sums_update_0_read_read_22_stage_127 <= dark_weights_weight_sums_update_0_read_read_22_stage_126;
      dark_weights_weight_sums_update_0_read_read_22_stage_128 <= dark_weights_weight_sums_update_0_read_read_22_stage_127;
      dark_weights_weight_sums_update_0_read_read_22_stage_129 <= dark_weights_weight_sums_update_0_read_read_22_stage_128;
      dark_weights_weight_sums_update_0_read_read_22_stage_130 <= dark_weights_weight_sums_update_0_read_read_22_stage_129;
      dark_weights_weight_sums_update_0_read_read_22_stage_131 <= dark_weights_weight_sums_update_0_read_read_22_stage_130;
      dark_weights_weight_sums_update_0_read_read_22_stage_132 <= dark_weights_weight_sums_update_0_read_read_22_stage_131;
      dark_weights_weight_sums_update_0_read_read_22_stage_133 <= dark_weights_weight_sums_update_0_read_read_22_stage_132;
      dark_weights_weight_sums_update_0_read_read_22_stage_134 <= dark_weights_weight_sums_update_0_read_read_22_stage_133;
      dark_weights_weight_sums_update_0_read_read_22_stage_135 <= dark_weights_weight_sums_update_0_read_read_22_stage_134;
      dark_weights_weight_sums_update_0_read_read_22_stage_136 <= dark_weights_weight_sums_update_0_read_read_22_stage_135;
      dark_weights_weight_sums_update_0_read_read_22_stage_137 <= dark_weights_weight_sums_update_0_read_read_22_stage_136;
      dark_weights_weight_sums_update_0_read_read_22_stage_138 <= dark_weights_weight_sums_update_0_read_read_22_stage_137;
      dark_weights_weight_sums_update_0_read_read_22_stage_139 <= dark_weights_weight_sums_update_0_read_read_22_stage_138;
      dark_weights_weight_sums_update_0_read_read_22_stage_140 <= dark_weights_weight_sums_update_0_read_read_22_stage_139;
      dark_weights_weight_sums_update_0_read_read_22_stage_141 <= dark_weights_weight_sums_update_0_read_read_22_stage_140;
      dark_weights_weight_sums_update_0_read_read_22_stage_142 <= dark_weights_weight_sums_update_0_read_read_22_stage_141;
      dark_weights_weight_sums_update_0_read_read_22_stage_143 <= dark_weights_weight_sums_update_0_read_read_22_stage_142;
      dark_weights_weight_sums_update_0_read_read_22_stage_144 <= dark_weights_weight_sums_update_0_read_read_22_stage_143;
      dark_weights_weight_sums_update_0_read_read_22_stage_145 <= dark_weights_weight_sums_update_0_read_read_22_stage_144;
      dark_weights_weight_sums_update_0_read_read_22_stage_146 <= dark_weights_weight_sums_update_0_read_read_22_stage_145;
      dark_weights_weight_sums_update_0_read_read_22_stage_147 <= dark_weights_weight_sums_update_0_read_read_22_stage_146;
      dark_weights_weight_sums_update_0_read_read_22_stage_148 <= dark_weights_weight_sums_update_0_read_read_22_stage_147;
      dark_weights_weight_sums_update_0_read_read_22_stage_149 <= dark_weights_weight_sums_update_0_read_read_22_stage_148;
      dark_weights_weight_sums_update_0_read_read_22_stage_150 <= dark_weights_weight_sums_update_0_read_read_22_stage_149;
      dark_weights_weight_sums_update_0_read_read_22_stage_151 <= dark_weights_weight_sums_update_0_read_read_22_stage_150;
      dark_weights_weight_sums_update_0_read_read_22_stage_152 <= dark_weights_weight_sums_update_0_read_read_22_stage_151;
      dark_weights_weight_sums_update_0_read_read_22_stage_153 <= dark_weights_weight_sums_update_0_read_read_22_stage_152;
      dark_weights_weight_sums_update_0_read_read_22_stage_154 <= dark_weights_weight_sums_update_0_read_read_22_stage_153;
      dark_weights_weight_sums_update_0_read_read_22_stage_155 <= dark_weights_weight_sums_update_0_read_read_22_stage_154;
      dark_weights_weight_sums_update_0_read_read_22_stage_156 <= dark_weights_weight_sums_update_0_read_read_22_stage_155;
      dark_weights_weight_sums_update_0_read_read_22_stage_157 <= dark_weights_weight_sums_update_0_read_read_22_stage_156;
      dark_weights_weight_sums_update_0_read_read_22_stage_158 <= dark_weights_weight_sums_update_0_read_read_22_stage_157;
      dark_weights_weight_sums_update_0_read_read_22_stage_159 <= dark_weights_weight_sums_update_0_read_read_22_stage_158;
      dark_weights_weight_sums_update_0_read_read_22_stage_160 <= dark_weights_weight_sums_update_0_read_read_22_stage_159;
      dark_weights_weight_sums_update_0_read_read_22_stage_161 <= dark_weights_weight_sums_update_0_read_read_22_stage_160;
      dark_weights_weight_sums_update_0_read_read_22_stage_162 <= dark_weights_weight_sums_update_0_read_read_22_stage_161;
      dark_weights_weight_sums_update_0_read_read_22_stage_163 <= dark_weights_weight_sums_update_0_read_read_22_stage_162;
      dark_weights_weight_sums_update_0_read_read_22_stage_164 <= dark_weights_weight_sums_update_0_read_read_22_stage_163;
      dark_weights_weight_sums_update_0_read_read_22_stage_165 <= dark_weights_weight_sums_update_0_read_read_22_stage_164;
      dark_weights_weight_sums_update_0_read_read_22_stage_166 <= dark_weights_weight_sums_update_0_read_read_22_stage_165;
      dark_weights_weight_sums_update_0_read_read_22_stage_167 <= dark_weights_weight_sums_update_0_read_read_22_stage_166;
      dark_weights_weight_sums_update_0_read_read_22_stage_168 <= dark_weights_weight_sums_update_0_read_read_22_stage_167;
      dark_weights_weight_sums_update_0_read_read_22_stage_169 <= dark_weights_weight_sums_update_0_read_read_22_stage_168;
      dark_weights_weight_sums_update_0_read_read_22_stage_170 <= dark_weights_weight_sums_update_0_read_read_22_stage_169;
      dark_weights_weight_sums_update_0_read_read_22_stage_171 <= dark_weights_weight_sums_update_0_read_read_22_stage_170;
      dark_weights_weight_sums_update_0_read_read_22_stage_172 <= dark_weights_weight_sums_update_0_read_read_22_stage_171;
      dark_weights_weight_sums_update_0_read_read_22_stage_173 <= dark_weights_weight_sums_update_0_read_read_22_stage_172;
      dark_weights_weight_sums_update_0_read_read_22_stage_174 <= dark_weights_weight_sums_update_0_read_read_22_stage_173;
      dark_weights_weight_sums_update_0_read_read_22_stage_175 <= dark_weights_weight_sums_update_0_read_read_22_stage_174;
      dark_weights_weight_sums_update_0_read_read_22_stage_176 <= dark_weights_weight_sums_update_0_read_read_22_stage_175;
      dark_weights_weight_sums_update_0_read_read_22_stage_177 <= dark_weights_weight_sums_update_0_read_read_22_stage_176;
      dark_weights_weight_sums_update_0_read_read_22_stage_178 <= dark_weights_weight_sums_update_0_read_read_22_stage_177;
      dark_weights_weight_sums_update_0_read_read_22_stage_179 <= dark_weights_weight_sums_update_0_read_read_22_stage_178;
      dark_weights_weight_sums_update_0_read_read_22_stage_180 <= dark_weights_weight_sums_update_0_read_read_22_stage_179;
      dark_weights_weight_sums_update_0_read_read_22_stage_181 <= dark_weights_weight_sums_update_0_read_read_22_stage_180;
      weight_sums_update_0_stage_37 <= weight_sums_update_0;
      weight_sums_update_0_stage_38 <= weight_sums_update_0_stage_37;
      weight_sums_update_0_stage_39 <= weight_sums_update_0_stage_38;
      weight_sums_update_0_stage_40 <= weight_sums_update_0_stage_39;
      weight_sums_update_0_stage_41 <= weight_sums_update_0_stage_40;
      weight_sums_update_0_stage_42 <= weight_sums_update_0_stage_41;
      weight_sums_update_0_stage_43 <= weight_sums_update_0_stage_42;
      weight_sums_update_0_stage_44 <= weight_sums_update_0_stage_43;
      weight_sums_update_0_stage_45 <= weight_sums_update_0_stage_44;
      weight_sums_update_0_stage_46 <= weight_sums_update_0_stage_45;
      weight_sums_update_0_stage_47 <= weight_sums_update_0_stage_46;
      weight_sums_update_0_stage_48 <= weight_sums_update_0_stage_47;
      weight_sums_update_0_stage_49 <= weight_sums_update_0_stage_48;
      weight_sums_update_0_stage_50 <= weight_sums_update_0_stage_49;
      weight_sums_update_0_stage_51 <= weight_sums_update_0_stage_50;
      weight_sums_update_0_stage_52 <= weight_sums_update_0_stage_51;
      weight_sums_update_0_stage_53 <= weight_sums_update_0_stage_52;
      weight_sums_update_0_stage_54 <= weight_sums_update_0_stage_53;
      weight_sums_update_0_stage_55 <= weight_sums_update_0_stage_54;
      weight_sums_update_0_stage_56 <= weight_sums_update_0_stage_55;
      weight_sums_update_0_stage_57 <= weight_sums_update_0_stage_56;
      weight_sums_update_0_stage_58 <= weight_sums_update_0_stage_57;
      weight_sums_update_0_stage_59 <= weight_sums_update_0_stage_58;
      weight_sums_update_0_stage_60 <= weight_sums_update_0_stage_59;
      weight_sums_update_0_stage_61 <= weight_sums_update_0_stage_60;
      weight_sums_update_0_stage_62 <= weight_sums_update_0_stage_61;
      weight_sums_update_0_stage_63 <= weight_sums_update_0_stage_62;
      weight_sums_update_0_stage_64 <= weight_sums_update_0_stage_63;
      weight_sums_update_0_stage_65 <= weight_sums_update_0_stage_64;
      weight_sums_update_0_stage_66 <= weight_sums_update_0_stage_65;
      weight_sums_update_0_stage_67 <= weight_sums_update_0_stage_66;
      weight_sums_update_0_stage_68 <= weight_sums_update_0_stage_67;
      weight_sums_update_0_stage_69 <= weight_sums_update_0_stage_68;
      weight_sums_update_0_stage_70 <= weight_sums_update_0_stage_69;
      weight_sums_update_0_stage_71 <= weight_sums_update_0_stage_70;
      weight_sums_update_0_stage_72 <= weight_sums_update_0_stage_71;
      weight_sums_update_0_stage_73 <= weight_sums_update_0_stage_72;
      weight_sums_update_0_stage_74 <= weight_sums_update_0_stage_73;
      weight_sums_update_0_stage_75 <= weight_sums_update_0_stage_74;
      weight_sums_update_0_stage_76 <= weight_sums_update_0_stage_75;
      weight_sums_update_0_stage_77 <= weight_sums_update_0_stage_76;
      weight_sums_update_0_stage_78 <= weight_sums_update_0_stage_77;
      weight_sums_update_0_stage_79 <= weight_sums_update_0_stage_78;
      weight_sums_update_0_stage_80 <= weight_sums_update_0_stage_79;
      weight_sums_update_0_stage_81 <= weight_sums_update_0_stage_80;
      weight_sums_update_0_stage_82 <= weight_sums_update_0_stage_81;
      weight_sums_update_0_stage_83 <= weight_sums_update_0_stage_82;
      weight_sums_update_0_stage_84 <= weight_sums_update_0_stage_83;
      weight_sums_update_0_stage_85 <= weight_sums_update_0_stage_84;
      weight_sums_update_0_stage_86 <= weight_sums_update_0_stage_85;
      weight_sums_update_0_stage_87 <= weight_sums_update_0_stage_86;
      weight_sums_update_0_stage_88 <= weight_sums_update_0_stage_87;
      weight_sums_update_0_stage_89 <= weight_sums_update_0_stage_88;
      weight_sums_update_0_stage_90 <= weight_sums_update_0_stage_89;
      weight_sums_update_0_stage_91 <= weight_sums_update_0_stage_90;
      weight_sums_update_0_stage_92 <= weight_sums_update_0_stage_91;
      weight_sums_update_0_stage_93 <= weight_sums_update_0_stage_92;
      weight_sums_update_0_stage_94 <= weight_sums_update_0_stage_93;
      weight_sums_update_0_stage_95 <= weight_sums_update_0_stage_94;
      weight_sums_update_0_stage_96 <= weight_sums_update_0_stage_95;
      weight_sums_update_0_stage_97 <= weight_sums_update_0_stage_96;
      weight_sums_update_0_stage_98 <= weight_sums_update_0_stage_97;
      weight_sums_update_0_stage_99 <= weight_sums_update_0_stage_98;
      weight_sums_update_0_stage_100 <= weight_sums_update_0_stage_99;
      weight_sums_update_0_stage_101 <= weight_sums_update_0_stage_100;
      weight_sums_update_0_stage_102 <= weight_sums_update_0_stage_101;
      weight_sums_update_0_stage_103 <= weight_sums_update_0_stage_102;
      weight_sums_update_0_stage_104 <= weight_sums_update_0_stage_103;
      weight_sums_update_0_stage_105 <= weight_sums_update_0_stage_104;
      weight_sums_update_0_stage_106 <= weight_sums_update_0_stage_105;
      weight_sums_update_0_stage_107 <= weight_sums_update_0_stage_106;
      weight_sums_update_0_stage_108 <= weight_sums_update_0_stage_107;
      weight_sums_update_0_stage_109 <= weight_sums_update_0_stage_108;
      weight_sums_update_0_stage_110 <= weight_sums_update_0_stage_109;
      weight_sums_update_0_stage_111 <= weight_sums_update_0_stage_110;
      weight_sums_update_0_stage_112 <= weight_sums_update_0_stage_111;
      weight_sums_update_0_stage_113 <= weight_sums_update_0_stage_112;
      weight_sums_update_0_stage_114 <= weight_sums_update_0_stage_113;
      weight_sums_update_0_stage_115 <= weight_sums_update_0_stage_114;
      weight_sums_update_0_stage_116 <= weight_sums_update_0_stage_115;
      weight_sums_update_0_stage_117 <= weight_sums_update_0_stage_116;
      weight_sums_update_0_stage_118 <= weight_sums_update_0_stage_117;
      weight_sums_update_0_stage_119 <= weight_sums_update_0_stage_118;
      weight_sums_update_0_stage_120 <= weight_sums_update_0_stage_119;
      weight_sums_update_0_stage_121 <= weight_sums_update_0_stage_120;
      weight_sums_update_0_stage_122 <= weight_sums_update_0_stage_121;
      weight_sums_update_0_stage_123 <= weight_sums_update_0_stage_122;
      weight_sums_update_0_stage_124 <= weight_sums_update_0_stage_123;
      weight_sums_update_0_stage_125 <= weight_sums_update_0_stage_124;
      weight_sums_update_0_stage_126 <= weight_sums_update_0_stage_125;
      weight_sums_update_0_stage_127 <= weight_sums_update_0_stage_126;
      weight_sums_update_0_stage_128 <= weight_sums_update_0_stage_127;
      weight_sums_update_0_stage_129 <= weight_sums_update_0_stage_128;
      weight_sums_update_0_stage_130 <= weight_sums_update_0_stage_129;
      weight_sums_update_0_stage_131 <= weight_sums_update_0_stage_130;
      weight_sums_update_0_stage_132 <= weight_sums_update_0_stage_131;
      weight_sums_update_0_stage_133 <= weight_sums_update_0_stage_132;
      weight_sums_update_0_stage_134 <= weight_sums_update_0_stage_133;
      weight_sums_update_0_stage_135 <= weight_sums_update_0_stage_134;
      weight_sums_update_0_stage_136 <= weight_sums_update_0_stage_135;
      weight_sums_update_0_stage_137 <= weight_sums_update_0_stage_136;
      weight_sums_update_0_stage_138 <= weight_sums_update_0_stage_137;
      weight_sums_update_0_stage_139 <= weight_sums_update_0_stage_138;
      weight_sums_update_0_stage_140 <= weight_sums_update_0_stage_139;
      weight_sums_update_0_stage_141 <= weight_sums_update_0_stage_140;
      weight_sums_update_0_stage_142 <= weight_sums_update_0_stage_141;
      weight_sums_update_0_stage_143 <= weight_sums_update_0_stage_142;
      weight_sums_update_0_stage_144 <= weight_sums_update_0_stage_143;
      weight_sums_update_0_stage_145 <= weight_sums_update_0_stage_144;
      weight_sums_update_0_stage_146 <= weight_sums_update_0_stage_145;
      weight_sums_update_0_stage_147 <= weight_sums_update_0_stage_146;
      weight_sums_update_0_stage_148 <= weight_sums_update_0_stage_147;
      weight_sums_update_0_stage_149 <= weight_sums_update_0_stage_148;
      weight_sums_update_0_stage_150 <= weight_sums_update_0_stage_149;
      weight_sums_update_0_stage_151 <= weight_sums_update_0_stage_150;
      weight_sums_update_0_stage_152 <= weight_sums_update_0_stage_151;
      weight_sums_update_0_stage_153 <= weight_sums_update_0_stage_152;
      weight_sums_update_0_stage_154 <= weight_sums_update_0_stage_153;
      weight_sums_update_0_stage_155 <= weight_sums_update_0_stage_154;
      weight_sums_update_0_stage_156 <= weight_sums_update_0_stage_155;
      weight_sums_update_0_stage_157 <= weight_sums_update_0_stage_156;
      weight_sums_update_0_stage_158 <= weight_sums_update_0_stage_157;
      weight_sums_update_0_stage_159 <= weight_sums_update_0_stage_158;
      weight_sums_update_0_stage_160 <= weight_sums_update_0_stage_159;
      weight_sums_update_0_stage_161 <= weight_sums_update_0_stage_160;
      weight_sums_update_0_stage_162 <= weight_sums_update_0_stage_161;
      weight_sums_update_0_stage_163 <= weight_sums_update_0_stage_162;
      weight_sums_update_0_stage_164 <= weight_sums_update_0_stage_163;
      weight_sums_update_0_stage_165 <= weight_sums_update_0_stage_164;
      weight_sums_update_0_stage_166 <= weight_sums_update_0_stage_165;
      weight_sums_update_0_stage_167 <= weight_sums_update_0_stage_166;
      weight_sums_update_0_stage_168 <= weight_sums_update_0_stage_167;
      weight_sums_update_0_stage_169 <= weight_sums_update_0_stage_168;
      weight_sums_update_0_stage_170 <= weight_sums_update_0_stage_169;
      weight_sums_update_0_stage_171 <= weight_sums_update_0_stage_170;
      weight_sums_update_0_stage_172 <= weight_sums_update_0_stage_171;
      weight_sums_update_0_stage_173 <= weight_sums_update_0_stage_172;
      weight_sums_update_0_stage_174 <= weight_sums_update_0_stage_173;
      weight_sums_update_0_stage_175 <= weight_sums_update_0_stage_174;
      weight_sums_update_0_stage_176 <= weight_sums_update_0_stage_175;
      weight_sums_update_0_stage_177 <= weight_sums_update_0_stage_176;
      weight_sums_update_0_stage_178 <= weight_sums_update_0_stage_177;
      weight_sums_update_0_stage_179 <= weight_sums_update_0_stage_178;
      weight_sums_update_0_stage_180 <= weight_sums_update_0_stage_179;
      weight_sums_update_0_stage_181 <= weight_sums_update_0_stage_180;
      bright_weights_weight_sums_update_0_read_read_23_stage_36 <= bright_weights_weight_sums_update_0_read_read_23;
      bright_weights_weight_sums_update_0_read_read_23_stage_37 <= bright_weights_weight_sums_update_0_read_read_23_stage_36;
      bright_weights_weight_sums_update_0_read_read_23_stage_38 <= bright_weights_weight_sums_update_0_read_read_23_stage_37;
      bright_weights_weight_sums_update_0_read_read_23_stage_39 <= bright_weights_weight_sums_update_0_read_read_23_stage_38;
      bright_weights_weight_sums_update_0_read_read_23_stage_40 <= bright_weights_weight_sums_update_0_read_read_23_stage_39;
      bright_weights_weight_sums_update_0_read_read_23_stage_41 <= bright_weights_weight_sums_update_0_read_read_23_stage_40;
      bright_weights_weight_sums_update_0_read_read_23_stage_42 <= bright_weights_weight_sums_update_0_read_read_23_stage_41;
      bright_weights_weight_sums_update_0_read_read_23_stage_43 <= bright_weights_weight_sums_update_0_read_read_23_stage_42;
      bright_weights_weight_sums_update_0_read_read_23_stage_44 <= bright_weights_weight_sums_update_0_read_read_23_stage_43;
      bright_weights_weight_sums_update_0_read_read_23_stage_45 <= bright_weights_weight_sums_update_0_read_read_23_stage_44;
      bright_weights_weight_sums_update_0_read_read_23_stage_46 <= bright_weights_weight_sums_update_0_read_read_23_stage_45;
      bright_weights_weight_sums_update_0_read_read_23_stage_47 <= bright_weights_weight_sums_update_0_read_read_23_stage_46;
      bright_weights_weight_sums_update_0_read_read_23_stage_48 <= bright_weights_weight_sums_update_0_read_read_23_stage_47;
      bright_weights_weight_sums_update_0_read_read_23_stage_49 <= bright_weights_weight_sums_update_0_read_read_23_stage_48;
      bright_weights_weight_sums_update_0_read_read_23_stage_50 <= bright_weights_weight_sums_update_0_read_read_23_stage_49;
      bright_weights_weight_sums_update_0_read_read_23_stage_51 <= bright_weights_weight_sums_update_0_read_read_23_stage_50;
      bright_weights_weight_sums_update_0_read_read_23_stage_52 <= bright_weights_weight_sums_update_0_read_read_23_stage_51;
      bright_weights_weight_sums_update_0_read_read_23_stage_53 <= bright_weights_weight_sums_update_0_read_read_23_stage_52;
      bright_weights_weight_sums_update_0_read_read_23_stage_54 <= bright_weights_weight_sums_update_0_read_read_23_stage_53;
      bright_weights_weight_sums_update_0_read_read_23_stage_55 <= bright_weights_weight_sums_update_0_read_read_23_stage_54;
      bright_weights_weight_sums_update_0_read_read_23_stage_56 <= bright_weights_weight_sums_update_0_read_read_23_stage_55;
      bright_weights_weight_sums_update_0_read_read_23_stage_57 <= bright_weights_weight_sums_update_0_read_read_23_stage_56;
      bright_weights_weight_sums_update_0_read_read_23_stage_58 <= bright_weights_weight_sums_update_0_read_read_23_stage_57;
      bright_weights_weight_sums_update_0_read_read_23_stage_59 <= bright_weights_weight_sums_update_0_read_read_23_stage_58;
      bright_weights_weight_sums_update_0_read_read_23_stage_60 <= bright_weights_weight_sums_update_0_read_read_23_stage_59;
      bright_weights_weight_sums_update_0_read_read_23_stage_61 <= bright_weights_weight_sums_update_0_read_read_23_stage_60;
      bright_weights_weight_sums_update_0_read_read_23_stage_62 <= bright_weights_weight_sums_update_0_read_read_23_stage_61;
      bright_weights_weight_sums_update_0_read_read_23_stage_63 <= bright_weights_weight_sums_update_0_read_read_23_stage_62;
      bright_weights_weight_sums_update_0_read_read_23_stage_64 <= bright_weights_weight_sums_update_0_read_read_23_stage_63;
      bright_weights_weight_sums_update_0_read_read_23_stage_65 <= bright_weights_weight_sums_update_0_read_read_23_stage_64;
      bright_weights_weight_sums_update_0_read_read_23_stage_66 <= bright_weights_weight_sums_update_0_read_read_23_stage_65;
      bright_weights_weight_sums_update_0_read_read_23_stage_67 <= bright_weights_weight_sums_update_0_read_read_23_stage_66;
      bright_weights_weight_sums_update_0_read_read_23_stage_68 <= bright_weights_weight_sums_update_0_read_read_23_stage_67;
      bright_weights_weight_sums_update_0_read_read_23_stage_69 <= bright_weights_weight_sums_update_0_read_read_23_stage_68;
      bright_weights_weight_sums_update_0_read_read_23_stage_70 <= bright_weights_weight_sums_update_0_read_read_23_stage_69;
      bright_weights_weight_sums_update_0_read_read_23_stage_71 <= bright_weights_weight_sums_update_0_read_read_23_stage_70;
      bright_weights_weight_sums_update_0_read_read_23_stage_72 <= bright_weights_weight_sums_update_0_read_read_23_stage_71;
      bright_weights_weight_sums_update_0_read_read_23_stage_73 <= bright_weights_weight_sums_update_0_read_read_23_stage_72;
      bright_weights_weight_sums_update_0_read_read_23_stage_74 <= bright_weights_weight_sums_update_0_read_read_23_stage_73;
      bright_weights_weight_sums_update_0_read_read_23_stage_75 <= bright_weights_weight_sums_update_0_read_read_23_stage_74;
      bright_weights_weight_sums_update_0_read_read_23_stage_76 <= bright_weights_weight_sums_update_0_read_read_23_stage_75;
      bright_weights_weight_sums_update_0_read_read_23_stage_77 <= bright_weights_weight_sums_update_0_read_read_23_stage_76;
      bright_weights_weight_sums_update_0_read_read_23_stage_78 <= bright_weights_weight_sums_update_0_read_read_23_stage_77;
      bright_weights_weight_sums_update_0_read_read_23_stage_79 <= bright_weights_weight_sums_update_0_read_read_23_stage_78;
      bright_weights_weight_sums_update_0_read_read_23_stage_80 <= bright_weights_weight_sums_update_0_read_read_23_stage_79;
      bright_weights_weight_sums_update_0_read_read_23_stage_81 <= bright_weights_weight_sums_update_0_read_read_23_stage_80;
      bright_weights_weight_sums_update_0_read_read_23_stage_82 <= bright_weights_weight_sums_update_0_read_read_23_stage_81;
      bright_weights_weight_sums_update_0_read_read_23_stage_83 <= bright_weights_weight_sums_update_0_read_read_23_stage_82;
      bright_weights_weight_sums_update_0_read_read_23_stage_84 <= bright_weights_weight_sums_update_0_read_read_23_stage_83;
      bright_weights_weight_sums_update_0_read_read_23_stage_85 <= bright_weights_weight_sums_update_0_read_read_23_stage_84;
      bright_weights_weight_sums_update_0_read_read_23_stage_86 <= bright_weights_weight_sums_update_0_read_read_23_stage_85;
      bright_weights_weight_sums_update_0_read_read_23_stage_87 <= bright_weights_weight_sums_update_0_read_read_23_stage_86;
      bright_weights_weight_sums_update_0_read_read_23_stage_88 <= bright_weights_weight_sums_update_0_read_read_23_stage_87;
      bright_weights_weight_sums_update_0_read_read_23_stage_89 <= bright_weights_weight_sums_update_0_read_read_23_stage_88;
      bright_weights_weight_sums_update_0_read_read_23_stage_90 <= bright_weights_weight_sums_update_0_read_read_23_stage_89;
      bright_weights_weight_sums_update_0_read_read_23_stage_91 <= bright_weights_weight_sums_update_0_read_read_23_stage_90;
      bright_weights_weight_sums_update_0_read_read_23_stage_92 <= bright_weights_weight_sums_update_0_read_read_23_stage_91;
      bright_weights_weight_sums_update_0_read_read_23_stage_93 <= bright_weights_weight_sums_update_0_read_read_23_stage_92;
      bright_weights_weight_sums_update_0_read_read_23_stage_94 <= bright_weights_weight_sums_update_0_read_read_23_stage_93;
      bright_weights_weight_sums_update_0_read_read_23_stage_95 <= bright_weights_weight_sums_update_0_read_read_23_stage_94;
      bright_weights_weight_sums_update_0_read_read_23_stage_96 <= bright_weights_weight_sums_update_0_read_read_23_stage_95;
      bright_weights_weight_sums_update_0_read_read_23_stage_97 <= bright_weights_weight_sums_update_0_read_read_23_stage_96;
      bright_weights_weight_sums_update_0_read_read_23_stage_98 <= bright_weights_weight_sums_update_0_read_read_23_stage_97;
      bright_weights_weight_sums_update_0_read_read_23_stage_99 <= bright_weights_weight_sums_update_0_read_read_23_stage_98;
      bright_weights_weight_sums_update_0_read_read_23_stage_100 <= bright_weights_weight_sums_update_0_read_read_23_stage_99;
      bright_weights_weight_sums_update_0_read_read_23_stage_101 <= bright_weights_weight_sums_update_0_read_read_23_stage_100;
      bright_weights_weight_sums_update_0_read_read_23_stage_102 <= bright_weights_weight_sums_update_0_read_read_23_stage_101;
      bright_weights_weight_sums_update_0_read_read_23_stage_103 <= bright_weights_weight_sums_update_0_read_read_23_stage_102;
      bright_weights_weight_sums_update_0_read_read_23_stage_104 <= bright_weights_weight_sums_update_0_read_read_23_stage_103;
      bright_weights_weight_sums_update_0_read_read_23_stage_105 <= bright_weights_weight_sums_update_0_read_read_23_stage_104;
      bright_weights_weight_sums_update_0_read_read_23_stage_106 <= bright_weights_weight_sums_update_0_read_read_23_stage_105;
      bright_weights_weight_sums_update_0_read_read_23_stage_107 <= bright_weights_weight_sums_update_0_read_read_23_stage_106;
      bright_weights_weight_sums_update_0_read_read_23_stage_108 <= bright_weights_weight_sums_update_0_read_read_23_stage_107;
      bright_weights_weight_sums_update_0_read_read_23_stage_109 <= bright_weights_weight_sums_update_0_read_read_23_stage_108;
      bright_weights_weight_sums_update_0_read_read_23_stage_110 <= bright_weights_weight_sums_update_0_read_read_23_stage_109;
      bright_weights_weight_sums_update_0_read_read_23_stage_111 <= bright_weights_weight_sums_update_0_read_read_23_stage_110;
      bright_weights_weight_sums_update_0_read_read_23_stage_112 <= bright_weights_weight_sums_update_0_read_read_23_stage_111;
      bright_weights_weight_sums_update_0_read_read_23_stage_113 <= bright_weights_weight_sums_update_0_read_read_23_stage_112;
      bright_weights_weight_sums_update_0_read_read_23_stage_114 <= bright_weights_weight_sums_update_0_read_read_23_stage_113;
      bright_weights_weight_sums_update_0_read_read_23_stage_115 <= bright_weights_weight_sums_update_0_read_read_23_stage_114;
      bright_weights_weight_sums_update_0_read_read_23_stage_116 <= bright_weights_weight_sums_update_0_read_read_23_stage_115;
      bright_weights_weight_sums_update_0_read_read_23_stage_117 <= bright_weights_weight_sums_update_0_read_read_23_stage_116;
      bright_weights_weight_sums_update_0_read_read_23_stage_118 <= bright_weights_weight_sums_update_0_read_read_23_stage_117;
      bright_weights_weight_sums_update_0_read_read_23_stage_119 <= bright_weights_weight_sums_update_0_read_read_23_stage_118;
      bright_weights_weight_sums_update_0_read_read_23_stage_120 <= bright_weights_weight_sums_update_0_read_read_23_stage_119;
      bright_weights_weight_sums_update_0_read_read_23_stage_121 <= bright_weights_weight_sums_update_0_read_read_23_stage_120;
      bright_weights_weight_sums_update_0_read_read_23_stage_122 <= bright_weights_weight_sums_update_0_read_read_23_stage_121;
      bright_weights_weight_sums_update_0_read_read_23_stage_123 <= bright_weights_weight_sums_update_0_read_read_23_stage_122;
      bright_weights_weight_sums_update_0_read_read_23_stage_124 <= bright_weights_weight_sums_update_0_read_read_23_stage_123;
      bright_weights_weight_sums_update_0_read_read_23_stage_125 <= bright_weights_weight_sums_update_0_read_read_23_stage_124;
      bright_weights_weight_sums_update_0_read_read_23_stage_126 <= bright_weights_weight_sums_update_0_read_read_23_stage_125;
      bright_weights_weight_sums_update_0_read_read_23_stage_127 <= bright_weights_weight_sums_update_0_read_read_23_stage_126;
      bright_weights_weight_sums_update_0_read_read_23_stage_128 <= bright_weights_weight_sums_update_0_read_read_23_stage_127;
      bright_weights_weight_sums_update_0_read_read_23_stage_129 <= bright_weights_weight_sums_update_0_read_read_23_stage_128;
      bright_weights_weight_sums_update_0_read_read_23_stage_130 <= bright_weights_weight_sums_update_0_read_read_23_stage_129;
      bright_weights_weight_sums_update_0_read_read_23_stage_131 <= bright_weights_weight_sums_update_0_read_read_23_stage_130;
      bright_weights_weight_sums_update_0_read_read_23_stage_132 <= bright_weights_weight_sums_update_0_read_read_23_stage_131;
      bright_weights_weight_sums_update_0_read_read_23_stage_133 <= bright_weights_weight_sums_update_0_read_read_23_stage_132;
      bright_weights_weight_sums_update_0_read_read_23_stage_134 <= bright_weights_weight_sums_update_0_read_read_23_stage_133;
      bright_weights_weight_sums_update_0_read_read_23_stage_135 <= bright_weights_weight_sums_update_0_read_read_23_stage_134;
      bright_weights_weight_sums_update_0_read_read_23_stage_136 <= bright_weights_weight_sums_update_0_read_read_23_stage_135;
      bright_weights_weight_sums_update_0_read_read_23_stage_137 <= bright_weights_weight_sums_update_0_read_read_23_stage_136;
      bright_weights_weight_sums_update_0_read_read_23_stage_138 <= bright_weights_weight_sums_update_0_read_read_23_stage_137;
      bright_weights_weight_sums_update_0_read_read_23_stage_139 <= bright_weights_weight_sums_update_0_read_read_23_stage_138;
      bright_weights_weight_sums_update_0_read_read_23_stage_140 <= bright_weights_weight_sums_update_0_read_read_23_stage_139;
      bright_weights_weight_sums_update_0_read_read_23_stage_141 <= bright_weights_weight_sums_update_0_read_read_23_stage_140;
      bright_weights_weight_sums_update_0_read_read_23_stage_142 <= bright_weights_weight_sums_update_0_read_read_23_stage_141;
      bright_weights_weight_sums_update_0_read_read_23_stage_143 <= bright_weights_weight_sums_update_0_read_read_23_stage_142;
      bright_weights_weight_sums_update_0_read_read_23_stage_144 <= bright_weights_weight_sums_update_0_read_read_23_stage_143;
      bright_weights_weight_sums_update_0_read_read_23_stage_145 <= bright_weights_weight_sums_update_0_read_read_23_stage_144;
      bright_weights_weight_sums_update_0_read_read_23_stage_146 <= bright_weights_weight_sums_update_0_read_read_23_stage_145;
      bright_weights_weight_sums_update_0_read_read_23_stage_147 <= bright_weights_weight_sums_update_0_read_read_23_stage_146;
      bright_weights_weight_sums_update_0_read_read_23_stage_148 <= bright_weights_weight_sums_update_0_read_read_23_stage_147;
      bright_weights_weight_sums_update_0_read_read_23_stage_149 <= bright_weights_weight_sums_update_0_read_read_23_stage_148;
      bright_weights_weight_sums_update_0_read_read_23_stage_150 <= bright_weights_weight_sums_update_0_read_read_23_stage_149;
      bright_weights_weight_sums_update_0_read_read_23_stage_151 <= bright_weights_weight_sums_update_0_read_read_23_stage_150;
      bright_weights_weight_sums_update_0_read_read_23_stage_152 <= bright_weights_weight_sums_update_0_read_read_23_stage_151;
      bright_weights_weight_sums_update_0_read_read_23_stage_153 <= bright_weights_weight_sums_update_0_read_read_23_stage_152;
      bright_weights_weight_sums_update_0_read_read_23_stage_154 <= bright_weights_weight_sums_update_0_read_read_23_stage_153;
      bright_weights_weight_sums_update_0_read_read_23_stage_155 <= bright_weights_weight_sums_update_0_read_read_23_stage_154;
      bright_weights_weight_sums_update_0_read_read_23_stage_156 <= bright_weights_weight_sums_update_0_read_read_23_stage_155;
      bright_weights_weight_sums_update_0_read_read_23_stage_157 <= bright_weights_weight_sums_update_0_read_read_23_stage_156;
      bright_weights_weight_sums_update_0_read_read_23_stage_158 <= bright_weights_weight_sums_update_0_read_read_23_stage_157;
      bright_weights_weight_sums_update_0_read_read_23_stage_159 <= bright_weights_weight_sums_update_0_read_read_23_stage_158;
      bright_weights_weight_sums_update_0_read_read_23_stage_160 <= bright_weights_weight_sums_update_0_read_read_23_stage_159;
      bright_weights_weight_sums_update_0_read_read_23_stage_161 <= bright_weights_weight_sums_update_0_read_read_23_stage_160;
      bright_weights_weight_sums_update_0_read_read_23_stage_162 <= bright_weights_weight_sums_update_0_read_read_23_stage_161;
      bright_weights_weight_sums_update_0_read_read_23_stage_163 <= bright_weights_weight_sums_update_0_read_read_23_stage_162;
      bright_weights_weight_sums_update_0_read_read_23_stage_164 <= bright_weights_weight_sums_update_0_read_read_23_stage_163;
      bright_weights_weight_sums_update_0_read_read_23_stage_165 <= bright_weights_weight_sums_update_0_read_read_23_stage_164;
      bright_weights_weight_sums_update_0_read_read_23_stage_166 <= bright_weights_weight_sums_update_0_read_read_23_stage_165;
      bright_weights_weight_sums_update_0_read_read_23_stage_167 <= bright_weights_weight_sums_update_0_read_read_23_stage_166;
      bright_weights_weight_sums_update_0_read_read_23_stage_168 <= bright_weights_weight_sums_update_0_read_read_23_stage_167;
      bright_weights_weight_sums_update_0_read_read_23_stage_169 <= bright_weights_weight_sums_update_0_read_read_23_stage_168;
      bright_weights_weight_sums_update_0_read_read_23_stage_170 <= bright_weights_weight_sums_update_0_read_read_23_stage_169;
      bright_weights_weight_sums_update_0_read_read_23_stage_171 <= bright_weights_weight_sums_update_0_read_read_23_stage_170;
      bright_weights_weight_sums_update_0_read_read_23_stage_172 <= bright_weights_weight_sums_update_0_read_read_23_stage_171;
      bright_weights_weight_sums_update_0_read_read_23_stage_173 <= bright_weights_weight_sums_update_0_read_read_23_stage_172;
      bright_weights_weight_sums_update_0_read_read_23_stage_174 <= bright_weights_weight_sums_update_0_read_read_23_stage_173;
      bright_weights_weight_sums_update_0_read_read_23_stage_175 <= bright_weights_weight_sums_update_0_read_read_23_stage_174;
      bright_weights_weight_sums_update_0_read_read_23_stage_176 <= bright_weights_weight_sums_update_0_read_read_23_stage_175;
      bright_weights_weight_sums_update_0_read_read_23_stage_177 <= bright_weights_weight_sums_update_0_read_read_23_stage_176;
      bright_weights_weight_sums_update_0_read_read_23_stage_178 <= bright_weights_weight_sums_update_0_read_read_23_stage_177;
      bright_weights_weight_sums_update_0_read_read_23_stage_179 <= bright_weights_weight_sums_update_0_read_read_23_stage_178;
      bright_weights_weight_sums_update_0_read_read_23_stage_180 <= bright_weights_weight_sums_update_0_read_read_23_stage_179;
      bright_weights_weight_sums_update_0_read_read_23_stage_181 <= bright_weights_weight_sums_update_0_read_read_23_stage_180;
      weight_sums_weight_sums_update_0_write_write_24_stage_38 <= weight_sums_weight_sums_update_0_write_write_24;
      weight_sums_weight_sums_update_0_write_write_24_stage_39 <= weight_sums_weight_sums_update_0_write_write_24_stage_38;
      weight_sums_weight_sums_update_0_write_write_24_stage_40 <= weight_sums_weight_sums_update_0_write_write_24_stage_39;
      weight_sums_weight_sums_update_0_write_write_24_stage_41 <= weight_sums_weight_sums_update_0_write_write_24_stage_40;
      weight_sums_weight_sums_update_0_write_write_24_stage_42 <= weight_sums_weight_sums_update_0_write_write_24_stage_41;
      weight_sums_weight_sums_update_0_write_write_24_stage_43 <= weight_sums_weight_sums_update_0_write_write_24_stage_42;
      weight_sums_weight_sums_update_0_write_write_24_stage_44 <= weight_sums_weight_sums_update_0_write_write_24_stage_43;
      weight_sums_weight_sums_update_0_write_write_24_stage_45 <= weight_sums_weight_sums_update_0_write_write_24_stage_44;
      weight_sums_weight_sums_update_0_write_write_24_stage_46 <= weight_sums_weight_sums_update_0_write_write_24_stage_45;
      weight_sums_weight_sums_update_0_write_write_24_stage_47 <= weight_sums_weight_sums_update_0_write_write_24_stage_46;
      weight_sums_weight_sums_update_0_write_write_24_stage_48 <= weight_sums_weight_sums_update_0_write_write_24_stage_47;
      weight_sums_weight_sums_update_0_write_write_24_stage_49 <= weight_sums_weight_sums_update_0_write_write_24_stage_48;
      weight_sums_weight_sums_update_0_write_write_24_stage_50 <= weight_sums_weight_sums_update_0_write_write_24_stage_49;
      weight_sums_weight_sums_update_0_write_write_24_stage_51 <= weight_sums_weight_sums_update_0_write_write_24_stage_50;
      weight_sums_weight_sums_update_0_write_write_24_stage_52 <= weight_sums_weight_sums_update_0_write_write_24_stage_51;
      weight_sums_weight_sums_update_0_write_write_24_stage_53 <= weight_sums_weight_sums_update_0_write_write_24_stage_52;
      weight_sums_weight_sums_update_0_write_write_24_stage_54 <= weight_sums_weight_sums_update_0_write_write_24_stage_53;
      weight_sums_weight_sums_update_0_write_write_24_stage_55 <= weight_sums_weight_sums_update_0_write_write_24_stage_54;
      weight_sums_weight_sums_update_0_write_write_24_stage_56 <= weight_sums_weight_sums_update_0_write_write_24_stage_55;
      weight_sums_weight_sums_update_0_write_write_24_stage_57 <= weight_sums_weight_sums_update_0_write_write_24_stage_56;
      weight_sums_weight_sums_update_0_write_write_24_stage_58 <= weight_sums_weight_sums_update_0_write_write_24_stage_57;
      weight_sums_weight_sums_update_0_write_write_24_stage_59 <= weight_sums_weight_sums_update_0_write_write_24_stage_58;
      weight_sums_weight_sums_update_0_write_write_24_stage_60 <= weight_sums_weight_sums_update_0_write_write_24_stage_59;
      weight_sums_weight_sums_update_0_write_write_24_stage_61 <= weight_sums_weight_sums_update_0_write_write_24_stage_60;
      weight_sums_weight_sums_update_0_write_write_24_stage_62 <= weight_sums_weight_sums_update_0_write_write_24_stage_61;
      weight_sums_weight_sums_update_0_write_write_24_stage_63 <= weight_sums_weight_sums_update_0_write_write_24_stage_62;
      weight_sums_weight_sums_update_0_write_write_24_stage_64 <= weight_sums_weight_sums_update_0_write_write_24_stage_63;
      weight_sums_weight_sums_update_0_write_write_24_stage_65 <= weight_sums_weight_sums_update_0_write_write_24_stage_64;
      weight_sums_weight_sums_update_0_write_write_24_stage_66 <= weight_sums_weight_sums_update_0_write_write_24_stage_65;
      weight_sums_weight_sums_update_0_write_write_24_stage_67 <= weight_sums_weight_sums_update_0_write_write_24_stage_66;
      weight_sums_weight_sums_update_0_write_write_24_stage_68 <= weight_sums_weight_sums_update_0_write_write_24_stage_67;
      weight_sums_weight_sums_update_0_write_write_24_stage_69 <= weight_sums_weight_sums_update_0_write_write_24_stage_68;
      weight_sums_weight_sums_update_0_write_write_24_stage_70 <= weight_sums_weight_sums_update_0_write_write_24_stage_69;
      weight_sums_weight_sums_update_0_write_write_24_stage_71 <= weight_sums_weight_sums_update_0_write_write_24_stage_70;
      weight_sums_weight_sums_update_0_write_write_24_stage_72 <= weight_sums_weight_sums_update_0_write_write_24_stage_71;
      weight_sums_weight_sums_update_0_write_write_24_stage_73 <= weight_sums_weight_sums_update_0_write_write_24_stage_72;
      weight_sums_weight_sums_update_0_write_write_24_stage_74 <= weight_sums_weight_sums_update_0_write_write_24_stage_73;
      weight_sums_weight_sums_update_0_write_write_24_stage_75 <= weight_sums_weight_sums_update_0_write_write_24_stage_74;
      weight_sums_weight_sums_update_0_write_write_24_stage_76 <= weight_sums_weight_sums_update_0_write_write_24_stage_75;
      weight_sums_weight_sums_update_0_write_write_24_stage_77 <= weight_sums_weight_sums_update_0_write_write_24_stage_76;
      weight_sums_weight_sums_update_0_write_write_24_stage_78 <= weight_sums_weight_sums_update_0_write_write_24_stage_77;
      weight_sums_weight_sums_update_0_write_write_24_stage_79 <= weight_sums_weight_sums_update_0_write_write_24_stage_78;
      weight_sums_weight_sums_update_0_write_write_24_stage_80 <= weight_sums_weight_sums_update_0_write_write_24_stage_79;
      weight_sums_weight_sums_update_0_write_write_24_stage_81 <= weight_sums_weight_sums_update_0_write_write_24_stage_80;
      weight_sums_weight_sums_update_0_write_write_24_stage_82 <= weight_sums_weight_sums_update_0_write_write_24_stage_81;
      weight_sums_weight_sums_update_0_write_write_24_stage_83 <= weight_sums_weight_sums_update_0_write_write_24_stage_82;
      weight_sums_weight_sums_update_0_write_write_24_stage_84 <= weight_sums_weight_sums_update_0_write_write_24_stage_83;
      weight_sums_weight_sums_update_0_write_write_24_stage_85 <= weight_sums_weight_sums_update_0_write_write_24_stage_84;
      weight_sums_weight_sums_update_0_write_write_24_stage_86 <= weight_sums_weight_sums_update_0_write_write_24_stage_85;
      weight_sums_weight_sums_update_0_write_write_24_stage_87 <= weight_sums_weight_sums_update_0_write_write_24_stage_86;
      weight_sums_weight_sums_update_0_write_write_24_stage_88 <= weight_sums_weight_sums_update_0_write_write_24_stage_87;
      weight_sums_weight_sums_update_0_write_write_24_stage_89 <= weight_sums_weight_sums_update_0_write_write_24_stage_88;
      weight_sums_weight_sums_update_0_write_write_24_stage_90 <= weight_sums_weight_sums_update_0_write_write_24_stage_89;
      weight_sums_weight_sums_update_0_write_write_24_stage_91 <= weight_sums_weight_sums_update_0_write_write_24_stage_90;
      weight_sums_weight_sums_update_0_write_write_24_stage_92 <= weight_sums_weight_sums_update_0_write_write_24_stage_91;
      weight_sums_weight_sums_update_0_write_write_24_stage_93 <= weight_sums_weight_sums_update_0_write_write_24_stage_92;
      weight_sums_weight_sums_update_0_write_write_24_stage_94 <= weight_sums_weight_sums_update_0_write_write_24_stage_93;
      weight_sums_weight_sums_update_0_write_write_24_stage_95 <= weight_sums_weight_sums_update_0_write_write_24_stage_94;
      weight_sums_weight_sums_update_0_write_write_24_stage_96 <= weight_sums_weight_sums_update_0_write_write_24_stage_95;
      weight_sums_weight_sums_update_0_write_write_24_stage_97 <= weight_sums_weight_sums_update_0_write_write_24_stage_96;
      weight_sums_weight_sums_update_0_write_write_24_stage_98 <= weight_sums_weight_sums_update_0_write_write_24_stage_97;
      weight_sums_weight_sums_update_0_write_write_24_stage_99 <= weight_sums_weight_sums_update_0_write_write_24_stage_98;
      weight_sums_weight_sums_update_0_write_write_24_stage_100 <= weight_sums_weight_sums_update_0_write_write_24_stage_99;
      weight_sums_weight_sums_update_0_write_write_24_stage_101 <= weight_sums_weight_sums_update_0_write_write_24_stage_100;
      weight_sums_weight_sums_update_0_write_write_24_stage_102 <= weight_sums_weight_sums_update_0_write_write_24_stage_101;
      weight_sums_weight_sums_update_0_write_write_24_stage_103 <= weight_sums_weight_sums_update_0_write_write_24_stage_102;
      weight_sums_weight_sums_update_0_write_write_24_stage_104 <= weight_sums_weight_sums_update_0_write_write_24_stage_103;
      weight_sums_weight_sums_update_0_write_write_24_stage_105 <= weight_sums_weight_sums_update_0_write_write_24_stage_104;
      weight_sums_weight_sums_update_0_write_write_24_stage_106 <= weight_sums_weight_sums_update_0_write_write_24_stage_105;
      weight_sums_weight_sums_update_0_write_write_24_stage_107 <= weight_sums_weight_sums_update_0_write_write_24_stage_106;
      weight_sums_weight_sums_update_0_write_write_24_stage_108 <= weight_sums_weight_sums_update_0_write_write_24_stage_107;
      weight_sums_weight_sums_update_0_write_write_24_stage_109 <= weight_sums_weight_sums_update_0_write_write_24_stage_108;
      weight_sums_weight_sums_update_0_write_write_24_stage_110 <= weight_sums_weight_sums_update_0_write_write_24_stage_109;
      weight_sums_weight_sums_update_0_write_write_24_stage_111 <= weight_sums_weight_sums_update_0_write_write_24_stage_110;
      weight_sums_weight_sums_update_0_write_write_24_stage_112 <= weight_sums_weight_sums_update_0_write_write_24_stage_111;
      weight_sums_weight_sums_update_0_write_write_24_stage_113 <= weight_sums_weight_sums_update_0_write_write_24_stage_112;
      weight_sums_weight_sums_update_0_write_write_24_stage_114 <= weight_sums_weight_sums_update_0_write_write_24_stage_113;
      weight_sums_weight_sums_update_0_write_write_24_stage_115 <= weight_sums_weight_sums_update_0_write_write_24_stage_114;
      weight_sums_weight_sums_update_0_write_write_24_stage_116 <= weight_sums_weight_sums_update_0_write_write_24_stage_115;
      weight_sums_weight_sums_update_0_write_write_24_stage_117 <= weight_sums_weight_sums_update_0_write_write_24_stage_116;
      weight_sums_weight_sums_update_0_write_write_24_stage_118 <= weight_sums_weight_sums_update_0_write_write_24_stage_117;
      weight_sums_weight_sums_update_0_write_write_24_stage_119 <= weight_sums_weight_sums_update_0_write_write_24_stage_118;
      weight_sums_weight_sums_update_0_write_write_24_stage_120 <= weight_sums_weight_sums_update_0_write_write_24_stage_119;
      weight_sums_weight_sums_update_0_write_write_24_stage_121 <= weight_sums_weight_sums_update_0_write_write_24_stage_120;
      weight_sums_weight_sums_update_0_write_write_24_stage_122 <= weight_sums_weight_sums_update_0_write_write_24_stage_121;
      weight_sums_weight_sums_update_0_write_write_24_stage_123 <= weight_sums_weight_sums_update_0_write_write_24_stage_122;
      weight_sums_weight_sums_update_0_write_write_24_stage_124 <= weight_sums_weight_sums_update_0_write_write_24_stage_123;
      weight_sums_weight_sums_update_0_write_write_24_stage_125 <= weight_sums_weight_sums_update_0_write_write_24_stage_124;
      weight_sums_weight_sums_update_0_write_write_24_stage_126 <= weight_sums_weight_sums_update_0_write_write_24_stage_125;
      weight_sums_weight_sums_update_0_write_write_24_stage_127 <= weight_sums_weight_sums_update_0_write_write_24_stage_126;
      weight_sums_weight_sums_update_0_write_write_24_stage_128 <= weight_sums_weight_sums_update_0_write_write_24_stage_127;
      weight_sums_weight_sums_update_0_write_write_24_stage_129 <= weight_sums_weight_sums_update_0_write_write_24_stage_128;
      weight_sums_weight_sums_update_0_write_write_24_stage_130 <= weight_sums_weight_sums_update_0_write_write_24_stage_129;
      weight_sums_weight_sums_update_0_write_write_24_stage_131 <= weight_sums_weight_sums_update_0_write_write_24_stage_130;
      weight_sums_weight_sums_update_0_write_write_24_stage_132 <= weight_sums_weight_sums_update_0_write_write_24_stage_131;
      weight_sums_weight_sums_update_0_write_write_24_stage_133 <= weight_sums_weight_sums_update_0_write_write_24_stage_132;
      weight_sums_weight_sums_update_0_write_write_24_stage_134 <= weight_sums_weight_sums_update_0_write_write_24_stage_133;
      weight_sums_weight_sums_update_0_write_write_24_stage_135 <= weight_sums_weight_sums_update_0_write_write_24_stage_134;
      weight_sums_weight_sums_update_0_write_write_24_stage_136 <= weight_sums_weight_sums_update_0_write_write_24_stage_135;
      weight_sums_weight_sums_update_0_write_write_24_stage_137 <= weight_sums_weight_sums_update_0_write_write_24_stage_136;
      weight_sums_weight_sums_update_0_write_write_24_stage_138 <= weight_sums_weight_sums_update_0_write_write_24_stage_137;
      weight_sums_weight_sums_update_0_write_write_24_stage_139 <= weight_sums_weight_sums_update_0_write_write_24_stage_138;
      weight_sums_weight_sums_update_0_write_write_24_stage_140 <= weight_sums_weight_sums_update_0_write_write_24_stage_139;
      weight_sums_weight_sums_update_0_write_write_24_stage_141 <= weight_sums_weight_sums_update_0_write_write_24_stage_140;
      weight_sums_weight_sums_update_0_write_write_24_stage_142 <= weight_sums_weight_sums_update_0_write_write_24_stage_141;
      weight_sums_weight_sums_update_0_write_write_24_stage_143 <= weight_sums_weight_sums_update_0_write_write_24_stage_142;
      weight_sums_weight_sums_update_0_write_write_24_stage_144 <= weight_sums_weight_sums_update_0_write_write_24_stage_143;
      weight_sums_weight_sums_update_0_write_write_24_stage_145 <= weight_sums_weight_sums_update_0_write_write_24_stage_144;
      weight_sums_weight_sums_update_0_write_write_24_stage_146 <= weight_sums_weight_sums_update_0_write_write_24_stage_145;
      weight_sums_weight_sums_update_0_write_write_24_stage_147 <= weight_sums_weight_sums_update_0_write_write_24_stage_146;
      weight_sums_weight_sums_update_0_write_write_24_stage_148 <= weight_sums_weight_sums_update_0_write_write_24_stage_147;
      weight_sums_weight_sums_update_0_write_write_24_stage_149 <= weight_sums_weight_sums_update_0_write_write_24_stage_148;
      weight_sums_weight_sums_update_0_write_write_24_stage_150 <= weight_sums_weight_sums_update_0_write_write_24_stage_149;
      weight_sums_weight_sums_update_0_write_write_24_stage_151 <= weight_sums_weight_sums_update_0_write_write_24_stage_150;
      weight_sums_weight_sums_update_0_write_write_24_stage_152 <= weight_sums_weight_sums_update_0_write_write_24_stage_151;
      weight_sums_weight_sums_update_0_write_write_24_stage_153 <= weight_sums_weight_sums_update_0_write_write_24_stage_152;
      weight_sums_weight_sums_update_0_write_write_24_stage_154 <= weight_sums_weight_sums_update_0_write_write_24_stage_153;
      weight_sums_weight_sums_update_0_write_write_24_stage_155 <= weight_sums_weight_sums_update_0_write_write_24_stage_154;
      weight_sums_weight_sums_update_0_write_write_24_stage_156 <= weight_sums_weight_sums_update_0_write_write_24_stage_155;
      weight_sums_weight_sums_update_0_write_write_24_stage_157 <= weight_sums_weight_sums_update_0_write_write_24_stage_156;
      weight_sums_weight_sums_update_0_write_write_24_stage_158 <= weight_sums_weight_sums_update_0_write_write_24_stage_157;
      weight_sums_weight_sums_update_0_write_write_24_stage_159 <= weight_sums_weight_sums_update_0_write_write_24_stage_158;
      weight_sums_weight_sums_update_0_write_write_24_stage_160 <= weight_sums_weight_sums_update_0_write_write_24_stage_159;
      weight_sums_weight_sums_update_0_write_write_24_stage_161 <= weight_sums_weight_sums_update_0_write_write_24_stage_160;
      weight_sums_weight_sums_update_0_write_write_24_stage_162 <= weight_sums_weight_sums_update_0_write_write_24_stage_161;
      weight_sums_weight_sums_update_0_write_write_24_stage_163 <= weight_sums_weight_sums_update_0_write_write_24_stage_162;
      weight_sums_weight_sums_update_0_write_write_24_stage_164 <= weight_sums_weight_sums_update_0_write_write_24_stage_163;
      weight_sums_weight_sums_update_0_write_write_24_stage_165 <= weight_sums_weight_sums_update_0_write_write_24_stage_164;
      weight_sums_weight_sums_update_0_write_write_24_stage_166 <= weight_sums_weight_sums_update_0_write_write_24_stage_165;
      weight_sums_weight_sums_update_0_write_write_24_stage_167 <= weight_sums_weight_sums_update_0_write_write_24_stage_166;
      weight_sums_weight_sums_update_0_write_write_24_stage_168 <= weight_sums_weight_sums_update_0_write_write_24_stage_167;
      weight_sums_weight_sums_update_0_write_write_24_stage_169 <= weight_sums_weight_sums_update_0_write_write_24_stage_168;
      weight_sums_weight_sums_update_0_write_write_24_stage_170 <= weight_sums_weight_sums_update_0_write_write_24_stage_169;
      weight_sums_weight_sums_update_0_write_write_24_stage_171 <= weight_sums_weight_sums_update_0_write_write_24_stage_170;
      weight_sums_weight_sums_update_0_write_write_24_stage_172 <= weight_sums_weight_sums_update_0_write_write_24_stage_171;
      weight_sums_weight_sums_update_0_write_write_24_stage_173 <= weight_sums_weight_sums_update_0_write_write_24_stage_172;
      weight_sums_weight_sums_update_0_write_write_24_stage_174 <= weight_sums_weight_sums_update_0_write_write_24_stage_173;
      weight_sums_weight_sums_update_0_write_write_24_stage_175 <= weight_sums_weight_sums_update_0_write_write_24_stage_174;
      weight_sums_weight_sums_update_0_write_write_24_stage_176 <= weight_sums_weight_sums_update_0_write_write_24_stage_175;
      weight_sums_weight_sums_update_0_write_write_24_stage_177 <= weight_sums_weight_sums_update_0_write_write_24_stage_176;
      weight_sums_weight_sums_update_0_write_write_24_stage_178 <= weight_sums_weight_sums_update_0_write_write_24_stage_177;
      weight_sums_weight_sums_update_0_write_write_24_stage_179 <= weight_sums_weight_sums_update_0_write_write_24_stage_178;
      weight_sums_weight_sums_update_0_write_write_24_stage_180 <= weight_sums_weight_sums_update_0_write_write_24_stage_179;
      weight_sums_weight_sums_update_0_write_write_24_stage_181 <= weight_sums_weight_sums_update_0_write_write_24_stage_180;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_42 <= dark_dark_laplace_diff_0_update_0_read_read_27;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_43 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_42;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_44 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_43;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_45 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_44;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_46 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_45;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_47 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_46;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_48 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_47;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_49 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_48;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_50 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_49;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_51 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_50;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_52 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_51;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_53 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_52;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_54 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_53;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_55 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_54;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_56 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_55;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_57 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_56;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_58 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_57;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_59 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_58;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_60 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_59;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_61 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_60;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_62 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_61;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_63 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_62;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_64 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_63;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_65 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_64;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_66 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_65;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_67 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_66;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_68 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_67;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_69 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_68;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_70 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_69;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_71 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_70;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_72 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_71;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_73 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_72;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_74 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_73;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_75 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_74;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_76 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_75;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_77 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_76;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_78 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_77;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_79 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_78;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_80 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_79;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_81 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_80;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_82 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_81;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_83 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_82;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_84 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_83;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_85 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_84;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_86 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_85;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_87 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_86;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_88 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_87;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_89 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_88;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_90 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_89;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_91 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_90;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_92 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_91;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_93 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_92;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_94 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_93;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_95 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_94;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_96 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_95;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_97 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_96;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_98 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_97;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_99 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_98;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_100 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_99;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_101 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_100;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_102 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_101;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_103 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_102;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_104 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_103;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_105 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_104;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_106 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_105;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_107 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_106;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_108 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_107;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_109 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_108;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_110 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_109;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_111 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_110;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_112 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_111;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_113 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_112;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_114 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_113;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_115 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_114;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_116 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_115;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_117 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_116;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_118 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_117;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_119 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_118;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_120 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_119;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_121 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_120;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_122 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_121;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_123 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_122;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_124 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_123;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_125 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_124;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_126 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_125;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_127 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_126;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_128 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_127;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_129 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_128;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_130 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_129;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_131 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_130;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_132 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_131;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_133 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_132;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_134 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_133;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_135 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_134;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_136 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_135;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_137 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_136;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_138 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_137;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_139 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_138;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_140 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_139;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_141 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_140;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_142 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_141;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_143 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_142;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_144 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_143;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_145 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_144;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_146 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_145;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_147 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_146;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_148 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_147;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_149 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_148;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_150 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_149;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_151 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_150;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_152 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_151;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_153 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_152;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_154 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_153;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_155 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_154;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_156 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_155;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_157 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_156;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_158 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_157;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_159 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_158;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_160 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_159;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_161 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_160;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_162 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_161;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_163 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_162;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_164 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_163;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_165 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_164;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_166 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_165;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_167 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_166;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_168 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_167;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_169 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_168;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_170 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_169;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_171 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_170;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_172 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_171;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_173 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_172;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_174 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_173;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_175 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_174;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_176 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_175;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_177 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_176;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_178 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_177;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_179 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_178;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_180 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_179;
      dark_dark_laplace_diff_0_update_0_read_read_27_stage_181 <= dark_dark_laplace_diff_0_update_0_read_read_27_stage_180;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_43 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_44 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_43;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_45 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_44;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_46 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_45;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_47 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_46;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_48 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_47;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_49 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_48;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_50 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_49;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_51 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_50;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_52 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_51;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_53 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_52;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_54 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_53;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_55 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_54;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_56 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_55;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_57 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_56;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_58 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_57;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_59 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_58;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_60 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_59;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_61 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_60;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_62 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_61;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_63 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_62;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_64 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_63;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_65 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_64;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_66 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_65;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_67 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_66;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_68 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_67;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_69 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_68;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_70 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_69;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_71 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_70;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_72 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_71;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_73 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_72;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_74 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_73;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_75 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_74;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_76 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_75;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_77 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_76;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_78 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_77;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_79 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_78;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_80 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_79;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_81 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_80;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_82 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_81;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_83 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_82;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_84 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_83;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_85 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_84;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_86 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_85;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_87 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_86;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_88 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_87;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_89 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_88;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_90 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_89;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_91 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_90;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_92 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_91;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_93 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_92;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_94 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_93;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_95 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_94;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_96 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_95;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_97 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_96;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_98 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_97;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_99 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_98;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_100 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_99;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_101 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_100;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_102 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_101;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_103 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_102;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_104 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_103;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_105 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_104;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_106 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_105;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_107 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_106;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_108 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_107;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_109 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_108;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_110 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_109;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_111 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_110;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_112 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_111;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_113 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_112;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_114 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_113;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_115 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_114;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_116 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_115;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_117 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_116;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_118 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_117;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_119 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_118;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_120 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_119;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_121 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_120;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_122 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_121;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_123 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_122;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_124 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_123;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_125 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_124;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_126 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_125;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_127 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_126;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_128 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_127;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_129 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_128;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_130 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_129;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_131 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_130;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_132 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_131;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_133 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_132;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_134 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_133;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_135 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_134;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_136 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_135;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_137 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_136;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_138 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_137;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_139 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_138;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_140 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_139;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_141 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_140;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_142 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_141;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_143 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_142;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_144 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_143;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_145 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_144;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_146 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_145;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_147 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_146;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_148 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_147;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_149 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_148;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_150 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_149;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_151 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_150;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_152 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_151;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_153 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_152;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_154 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_153;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_155 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_154;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_156 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_155;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_157 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_156;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_158 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_157;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_159 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_158;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_160 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_159;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_161 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_160;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_162 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_161;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_163 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_162;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_164 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_163;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_165 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_164;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_166 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_165;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_167 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_166;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_168 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_167;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_169 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_168;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_170 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_169;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_171 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_170;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_172 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_171;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_173 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_172;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_174 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_173;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_175 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_174;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_176 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_175;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_177 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_176;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_178 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_177;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_179 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_178;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_180 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_179;
      dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_181 <= dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28_stage_180;
      dark_laplace_diff_0_update_0_stage_44 <= dark_laplace_diff_0_update_0;
      dark_laplace_diff_0_update_0_stage_45 <= dark_laplace_diff_0_update_0_stage_44;
      dark_laplace_diff_0_update_0_stage_46 <= dark_laplace_diff_0_update_0_stage_45;
      dark_laplace_diff_0_update_0_stage_47 <= dark_laplace_diff_0_update_0_stage_46;
      dark_laplace_diff_0_update_0_stage_48 <= dark_laplace_diff_0_update_0_stage_47;
      dark_laplace_diff_0_update_0_stage_49 <= dark_laplace_diff_0_update_0_stage_48;
      dark_laplace_diff_0_update_0_stage_50 <= dark_laplace_diff_0_update_0_stage_49;
      dark_laplace_diff_0_update_0_stage_51 <= dark_laplace_diff_0_update_0_stage_50;
      dark_laplace_diff_0_update_0_stage_52 <= dark_laplace_diff_0_update_0_stage_51;
      dark_laplace_diff_0_update_0_stage_53 <= dark_laplace_diff_0_update_0_stage_52;
      dark_laplace_diff_0_update_0_stage_54 <= dark_laplace_diff_0_update_0_stage_53;
      dark_laplace_diff_0_update_0_stage_55 <= dark_laplace_diff_0_update_0_stage_54;
      dark_laplace_diff_0_update_0_stage_56 <= dark_laplace_diff_0_update_0_stage_55;
      dark_laplace_diff_0_update_0_stage_57 <= dark_laplace_diff_0_update_0_stage_56;
      dark_laplace_diff_0_update_0_stage_58 <= dark_laplace_diff_0_update_0_stage_57;
      dark_laplace_diff_0_update_0_stage_59 <= dark_laplace_diff_0_update_0_stage_58;
      dark_laplace_diff_0_update_0_stage_60 <= dark_laplace_diff_0_update_0_stage_59;
      dark_laplace_diff_0_update_0_stage_61 <= dark_laplace_diff_0_update_0_stage_60;
      dark_laplace_diff_0_update_0_stage_62 <= dark_laplace_diff_0_update_0_stage_61;
      dark_laplace_diff_0_update_0_stage_63 <= dark_laplace_diff_0_update_0_stage_62;
      dark_laplace_diff_0_update_0_stage_64 <= dark_laplace_diff_0_update_0_stage_63;
      dark_laplace_diff_0_update_0_stage_65 <= dark_laplace_diff_0_update_0_stage_64;
      dark_laplace_diff_0_update_0_stage_66 <= dark_laplace_diff_0_update_0_stage_65;
      dark_laplace_diff_0_update_0_stage_67 <= dark_laplace_diff_0_update_0_stage_66;
      dark_laplace_diff_0_update_0_stage_68 <= dark_laplace_diff_0_update_0_stage_67;
      dark_laplace_diff_0_update_0_stage_69 <= dark_laplace_diff_0_update_0_stage_68;
      dark_laplace_diff_0_update_0_stage_70 <= dark_laplace_diff_0_update_0_stage_69;
      dark_laplace_diff_0_update_0_stage_71 <= dark_laplace_diff_0_update_0_stage_70;
      dark_laplace_diff_0_update_0_stage_72 <= dark_laplace_diff_0_update_0_stage_71;
      dark_laplace_diff_0_update_0_stage_73 <= dark_laplace_diff_0_update_0_stage_72;
      dark_laplace_diff_0_update_0_stage_74 <= dark_laplace_diff_0_update_0_stage_73;
      dark_laplace_diff_0_update_0_stage_75 <= dark_laplace_diff_0_update_0_stage_74;
      dark_laplace_diff_0_update_0_stage_76 <= dark_laplace_diff_0_update_0_stage_75;
      dark_laplace_diff_0_update_0_stage_77 <= dark_laplace_diff_0_update_0_stage_76;
      dark_laplace_diff_0_update_0_stage_78 <= dark_laplace_diff_0_update_0_stage_77;
      dark_laplace_diff_0_update_0_stage_79 <= dark_laplace_diff_0_update_0_stage_78;
      dark_laplace_diff_0_update_0_stage_80 <= dark_laplace_diff_0_update_0_stage_79;
      dark_laplace_diff_0_update_0_stage_81 <= dark_laplace_diff_0_update_0_stage_80;
      dark_laplace_diff_0_update_0_stage_82 <= dark_laplace_diff_0_update_0_stage_81;
      dark_laplace_diff_0_update_0_stage_83 <= dark_laplace_diff_0_update_0_stage_82;
      dark_laplace_diff_0_update_0_stage_84 <= dark_laplace_diff_0_update_0_stage_83;
      dark_laplace_diff_0_update_0_stage_85 <= dark_laplace_diff_0_update_0_stage_84;
      dark_laplace_diff_0_update_0_stage_86 <= dark_laplace_diff_0_update_0_stage_85;
      dark_laplace_diff_0_update_0_stage_87 <= dark_laplace_diff_0_update_0_stage_86;
      dark_laplace_diff_0_update_0_stage_88 <= dark_laplace_diff_0_update_0_stage_87;
      dark_laplace_diff_0_update_0_stage_89 <= dark_laplace_diff_0_update_0_stage_88;
      dark_laplace_diff_0_update_0_stage_90 <= dark_laplace_diff_0_update_0_stage_89;
      dark_laplace_diff_0_update_0_stage_91 <= dark_laplace_diff_0_update_0_stage_90;
      dark_laplace_diff_0_update_0_stage_92 <= dark_laplace_diff_0_update_0_stage_91;
      dark_laplace_diff_0_update_0_stage_93 <= dark_laplace_diff_0_update_0_stage_92;
      dark_laplace_diff_0_update_0_stage_94 <= dark_laplace_diff_0_update_0_stage_93;
      dark_laplace_diff_0_update_0_stage_95 <= dark_laplace_diff_0_update_0_stage_94;
      dark_laplace_diff_0_update_0_stage_96 <= dark_laplace_diff_0_update_0_stage_95;
      dark_laplace_diff_0_update_0_stage_97 <= dark_laplace_diff_0_update_0_stage_96;
      dark_laplace_diff_0_update_0_stage_98 <= dark_laplace_diff_0_update_0_stage_97;
      dark_laplace_diff_0_update_0_stage_99 <= dark_laplace_diff_0_update_0_stage_98;
      dark_laplace_diff_0_update_0_stage_100 <= dark_laplace_diff_0_update_0_stage_99;
      dark_laplace_diff_0_update_0_stage_101 <= dark_laplace_diff_0_update_0_stage_100;
      dark_laplace_diff_0_update_0_stage_102 <= dark_laplace_diff_0_update_0_stage_101;
      dark_laplace_diff_0_update_0_stage_103 <= dark_laplace_diff_0_update_0_stage_102;
      dark_laplace_diff_0_update_0_stage_104 <= dark_laplace_diff_0_update_0_stage_103;
      dark_laplace_diff_0_update_0_stage_105 <= dark_laplace_diff_0_update_0_stage_104;
      dark_laplace_diff_0_update_0_stage_106 <= dark_laplace_diff_0_update_0_stage_105;
      dark_laplace_diff_0_update_0_stage_107 <= dark_laplace_diff_0_update_0_stage_106;
      dark_laplace_diff_0_update_0_stage_108 <= dark_laplace_diff_0_update_0_stage_107;
      dark_laplace_diff_0_update_0_stage_109 <= dark_laplace_diff_0_update_0_stage_108;
      dark_laplace_diff_0_update_0_stage_110 <= dark_laplace_diff_0_update_0_stage_109;
      dark_laplace_diff_0_update_0_stage_111 <= dark_laplace_diff_0_update_0_stage_110;
      dark_laplace_diff_0_update_0_stage_112 <= dark_laplace_diff_0_update_0_stage_111;
      dark_laplace_diff_0_update_0_stage_113 <= dark_laplace_diff_0_update_0_stage_112;
      dark_laplace_diff_0_update_0_stage_114 <= dark_laplace_diff_0_update_0_stage_113;
      dark_laplace_diff_0_update_0_stage_115 <= dark_laplace_diff_0_update_0_stage_114;
      dark_laplace_diff_0_update_0_stage_116 <= dark_laplace_diff_0_update_0_stage_115;
      dark_laplace_diff_0_update_0_stage_117 <= dark_laplace_diff_0_update_0_stage_116;
      dark_laplace_diff_0_update_0_stage_118 <= dark_laplace_diff_0_update_0_stage_117;
      dark_laplace_diff_0_update_0_stage_119 <= dark_laplace_diff_0_update_0_stage_118;
      dark_laplace_diff_0_update_0_stage_120 <= dark_laplace_diff_0_update_0_stage_119;
      dark_laplace_diff_0_update_0_stage_121 <= dark_laplace_diff_0_update_0_stage_120;
      dark_laplace_diff_0_update_0_stage_122 <= dark_laplace_diff_0_update_0_stage_121;
      dark_laplace_diff_0_update_0_stage_123 <= dark_laplace_diff_0_update_0_stage_122;
      dark_laplace_diff_0_update_0_stage_124 <= dark_laplace_diff_0_update_0_stage_123;
      dark_laplace_diff_0_update_0_stage_125 <= dark_laplace_diff_0_update_0_stage_124;
      dark_laplace_diff_0_update_0_stage_126 <= dark_laplace_diff_0_update_0_stage_125;
      dark_laplace_diff_0_update_0_stage_127 <= dark_laplace_diff_0_update_0_stage_126;
      dark_laplace_diff_0_update_0_stage_128 <= dark_laplace_diff_0_update_0_stage_127;
      dark_laplace_diff_0_update_0_stage_129 <= dark_laplace_diff_0_update_0_stage_128;
      dark_laplace_diff_0_update_0_stage_130 <= dark_laplace_diff_0_update_0_stage_129;
      dark_laplace_diff_0_update_0_stage_131 <= dark_laplace_diff_0_update_0_stage_130;
      dark_laplace_diff_0_update_0_stage_132 <= dark_laplace_diff_0_update_0_stage_131;
      dark_laplace_diff_0_update_0_stage_133 <= dark_laplace_diff_0_update_0_stage_132;
      dark_laplace_diff_0_update_0_stage_134 <= dark_laplace_diff_0_update_0_stage_133;
      dark_laplace_diff_0_update_0_stage_135 <= dark_laplace_diff_0_update_0_stage_134;
      dark_laplace_diff_0_update_0_stage_136 <= dark_laplace_diff_0_update_0_stage_135;
      dark_laplace_diff_0_update_0_stage_137 <= dark_laplace_diff_0_update_0_stage_136;
      dark_laplace_diff_0_update_0_stage_138 <= dark_laplace_diff_0_update_0_stage_137;
      dark_laplace_diff_0_update_0_stage_139 <= dark_laplace_diff_0_update_0_stage_138;
      dark_laplace_diff_0_update_0_stage_140 <= dark_laplace_diff_0_update_0_stage_139;
      dark_laplace_diff_0_update_0_stage_141 <= dark_laplace_diff_0_update_0_stage_140;
      dark_laplace_diff_0_update_0_stage_142 <= dark_laplace_diff_0_update_0_stage_141;
      dark_laplace_diff_0_update_0_stage_143 <= dark_laplace_diff_0_update_0_stage_142;
      dark_laplace_diff_0_update_0_stage_144 <= dark_laplace_diff_0_update_0_stage_143;
      dark_laplace_diff_0_update_0_stage_145 <= dark_laplace_diff_0_update_0_stage_144;
      dark_laplace_diff_0_update_0_stage_146 <= dark_laplace_diff_0_update_0_stage_145;
      dark_laplace_diff_0_update_0_stage_147 <= dark_laplace_diff_0_update_0_stage_146;
      dark_laplace_diff_0_update_0_stage_148 <= dark_laplace_diff_0_update_0_stage_147;
      dark_laplace_diff_0_update_0_stage_149 <= dark_laplace_diff_0_update_0_stage_148;
      dark_laplace_diff_0_update_0_stage_150 <= dark_laplace_diff_0_update_0_stage_149;
      dark_laplace_diff_0_update_0_stage_151 <= dark_laplace_diff_0_update_0_stage_150;
      dark_laplace_diff_0_update_0_stage_152 <= dark_laplace_diff_0_update_0_stage_151;
      dark_laplace_diff_0_update_0_stage_153 <= dark_laplace_diff_0_update_0_stage_152;
      dark_laplace_diff_0_update_0_stage_154 <= dark_laplace_diff_0_update_0_stage_153;
      dark_laplace_diff_0_update_0_stage_155 <= dark_laplace_diff_0_update_0_stage_154;
      dark_laplace_diff_0_update_0_stage_156 <= dark_laplace_diff_0_update_0_stage_155;
      dark_laplace_diff_0_update_0_stage_157 <= dark_laplace_diff_0_update_0_stage_156;
      dark_laplace_diff_0_update_0_stage_158 <= dark_laplace_diff_0_update_0_stage_157;
      dark_laplace_diff_0_update_0_stage_159 <= dark_laplace_diff_0_update_0_stage_158;
      dark_laplace_diff_0_update_0_stage_160 <= dark_laplace_diff_0_update_0_stage_159;
      dark_laplace_diff_0_update_0_stage_161 <= dark_laplace_diff_0_update_0_stage_160;
      dark_laplace_diff_0_update_0_stage_162 <= dark_laplace_diff_0_update_0_stage_161;
      dark_laplace_diff_0_update_0_stage_163 <= dark_laplace_diff_0_update_0_stage_162;
      dark_laplace_diff_0_update_0_stage_164 <= dark_laplace_diff_0_update_0_stage_163;
      dark_laplace_diff_0_update_0_stage_165 <= dark_laplace_diff_0_update_0_stage_164;
      dark_laplace_diff_0_update_0_stage_166 <= dark_laplace_diff_0_update_0_stage_165;
      dark_laplace_diff_0_update_0_stage_167 <= dark_laplace_diff_0_update_0_stage_166;
      dark_laplace_diff_0_update_0_stage_168 <= dark_laplace_diff_0_update_0_stage_167;
      dark_laplace_diff_0_update_0_stage_169 <= dark_laplace_diff_0_update_0_stage_168;
      dark_laplace_diff_0_update_0_stage_170 <= dark_laplace_diff_0_update_0_stage_169;
      dark_laplace_diff_0_update_0_stage_171 <= dark_laplace_diff_0_update_0_stage_170;
      dark_laplace_diff_0_update_0_stage_172 <= dark_laplace_diff_0_update_0_stage_171;
      dark_laplace_diff_0_update_0_stage_173 <= dark_laplace_diff_0_update_0_stage_172;
      dark_laplace_diff_0_update_0_stage_174 <= dark_laplace_diff_0_update_0_stage_173;
      dark_laplace_diff_0_update_0_stage_175 <= dark_laplace_diff_0_update_0_stage_174;
      dark_laplace_diff_0_update_0_stage_176 <= dark_laplace_diff_0_update_0_stage_175;
      dark_laplace_diff_0_update_0_stage_177 <= dark_laplace_diff_0_update_0_stage_176;
      dark_laplace_diff_0_update_0_stage_178 <= dark_laplace_diff_0_update_0_stage_177;
      dark_laplace_diff_0_update_0_stage_179 <= dark_laplace_diff_0_update_0_stage_178;
      dark_laplace_diff_0_update_0_stage_180 <= dark_laplace_diff_0_update_0_stage_179;
      dark_laplace_diff_0_update_0_stage_181 <= dark_laplace_diff_0_update_0_stage_180;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_45 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_46 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_45;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_47 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_46;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_48 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_47;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_49 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_48;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_50 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_49;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_51 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_50;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_52 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_51;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_53 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_52;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_54 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_53;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_55 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_54;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_56 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_55;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_57 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_56;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_58 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_57;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_59 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_58;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_60 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_59;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_61 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_60;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_62 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_61;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_63 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_62;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_64 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_63;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_65 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_64;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_66 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_65;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_67 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_66;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_68 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_67;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_69 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_68;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_70 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_69;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_71 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_70;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_72 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_71;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_73 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_72;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_74 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_73;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_75 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_74;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_76 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_75;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_77 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_76;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_78 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_77;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_79 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_78;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_80 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_79;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_81 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_80;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_82 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_81;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_83 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_82;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_84 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_83;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_85 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_84;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_86 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_85;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_87 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_86;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_88 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_87;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_89 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_88;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_90 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_89;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_91 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_90;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_92 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_91;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_93 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_92;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_94 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_93;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_95 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_94;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_96 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_95;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_97 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_96;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_98 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_97;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_99 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_98;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_100 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_99;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_101 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_100;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_102 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_101;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_103 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_102;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_104 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_103;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_105 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_104;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_106 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_105;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_107 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_106;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_108 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_107;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_109 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_108;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_110 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_109;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_111 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_110;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_112 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_111;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_113 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_112;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_114 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_113;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_115 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_114;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_116 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_115;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_117 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_116;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_118 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_117;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_119 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_118;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_120 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_119;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_121 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_120;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_122 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_121;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_123 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_122;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_124 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_123;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_125 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_124;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_126 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_125;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_127 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_126;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_128 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_127;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_129 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_128;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_130 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_129;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_131 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_130;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_132 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_131;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_133 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_132;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_134 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_133;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_135 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_134;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_136 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_135;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_137 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_136;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_138 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_137;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_139 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_138;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_140 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_139;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_141 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_140;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_142 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_141;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_143 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_142;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_144 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_143;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_145 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_144;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_146 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_145;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_147 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_146;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_148 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_147;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_149 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_148;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_150 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_149;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_151 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_150;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_152 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_151;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_153 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_152;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_154 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_153;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_155 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_154;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_156 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_155;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_157 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_156;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_158 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_157;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_159 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_158;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_160 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_159;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_161 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_160;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_162 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_161;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_163 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_162;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_164 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_163;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_165 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_164;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_166 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_165;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_167 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_166;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_168 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_167;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_169 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_168;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_170 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_169;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_171 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_170;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_172 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_171;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_173 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_172;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_174 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_173;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_175 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_174;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_176 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_175;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_177 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_176;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_178 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_177;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_179 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_178;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_180 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_179;
      dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_181 <= dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29_stage_180;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_49 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_50 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_49;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_51 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_50;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_52 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_51;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_53 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_52;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_54 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_53;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_55 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_54;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_56 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_55;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_57 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_56;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_58 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_57;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_59 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_58;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_60 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_59;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_61 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_60;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_62 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_61;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_63 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_62;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_64 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_63;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_65 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_64;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_66 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_65;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_67 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_66;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_68 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_67;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_69 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_68;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_70 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_69;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_71 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_70;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_72 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_71;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_73 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_72;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_74 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_73;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_75 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_74;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_76 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_75;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_77 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_76;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_78 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_77;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_79 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_78;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_80 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_79;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_81 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_80;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_82 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_81;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_83 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_82;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_84 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_83;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_85 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_84;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_86 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_85;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_87 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_86;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_88 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_87;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_89 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_88;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_90 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_89;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_91 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_90;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_92 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_91;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_93 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_92;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_94 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_93;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_95 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_94;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_96 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_95;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_97 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_96;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_98 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_97;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_99 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_98;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_100 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_99;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_101 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_100;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_102 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_101;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_103 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_102;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_104 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_103;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_105 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_104;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_106 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_105;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_107 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_106;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_108 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_107;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_109 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_108;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_110 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_109;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_111 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_110;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_112 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_111;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_113 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_112;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_114 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_113;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_115 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_114;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_116 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_115;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_117 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_116;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_118 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_117;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_119 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_118;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_120 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_119;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_121 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_120;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_122 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_121;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_123 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_122;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_124 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_123;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_125 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_124;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_126 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_125;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_127 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_126;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_128 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_127;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_129 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_128;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_130 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_129;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_131 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_130;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_132 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_131;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_133 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_132;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_134 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_133;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_135 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_134;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_136 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_135;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_137 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_136;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_138 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_137;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_139 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_138;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_140 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_139;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_141 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_140;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_142 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_141;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_143 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_142;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_144 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_143;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_145 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_144;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_146 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_145;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_147 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_146;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_148 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_147;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_149 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_148;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_150 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_149;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_151 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_150;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_152 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_151;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_153 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_152;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_154 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_153;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_155 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_154;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_156 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_155;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_157 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_156;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_158 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_157;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_159 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_158;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_160 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_159;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_161 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_160;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_162 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_161;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_163 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_162;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_164 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_163;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_165 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_164;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_166 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_165;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_167 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_166;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_168 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_167;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_169 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_168;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_170 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_169;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_171 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_170;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_172 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_171;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_173 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_172;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_174 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_173;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_175 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_174;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_176 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_175;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_177 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_176;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_178 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_177;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_179 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_178;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_180 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_179;
      bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_181 <= bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32_stage_180;
      bright_gauss_ds_2_update_0_stage_50 <= bright_gauss_ds_2_update_0;
      bright_gauss_ds_2_update_0_stage_51 <= bright_gauss_ds_2_update_0_stage_50;
      bright_gauss_ds_2_update_0_stage_52 <= bright_gauss_ds_2_update_0_stage_51;
      bright_gauss_ds_2_update_0_stage_53 <= bright_gauss_ds_2_update_0_stage_52;
      bright_gauss_ds_2_update_0_stage_54 <= bright_gauss_ds_2_update_0_stage_53;
      bright_gauss_ds_2_update_0_stage_55 <= bright_gauss_ds_2_update_0_stage_54;
      bright_gauss_ds_2_update_0_stage_56 <= bright_gauss_ds_2_update_0_stage_55;
      bright_gauss_ds_2_update_0_stage_57 <= bright_gauss_ds_2_update_0_stage_56;
      bright_gauss_ds_2_update_0_stage_58 <= bright_gauss_ds_2_update_0_stage_57;
      bright_gauss_ds_2_update_0_stage_59 <= bright_gauss_ds_2_update_0_stage_58;
      bright_gauss_ds_2_update_0_stage_60 <= bright_gauss_ds_2_update_0_stage_59;
      bright_gauss_ds_2_update_0_stage_61 <= bright_gauss_ds_2_update_0_stage_60;
      bright_gauss_ds_2_update_0_stage_62 <= bright_gauss_ds_2_update_0_stage_61;
      bright_gauss_ds_2_update_0_stage_63 <= bright_gauss_ds_2_update_0_stage_62;
      bright_gauss_ds_2_update_0_stage_64 <= bright_gauss_ds_2_update_0_stage_63;
      bright_gauss_ds_2_update_0_stage_65 <= bright_gauss_ds_2_update_0_stage_64;
      bright_gauss_ds_2_update_0_stage_66 <= bright_gauss_ds_2_update_0_stage_65;
      bright_gauss_ds_2_update_0_stage_67 <= bright_gauss_ds_2_update_0_stage_66;
      bright_gauss_ds_2_update_0_stage_68 <= bright_gauss_ds_2_update_0_stage_67;
      bright_gauss_ds_2_update_0_stage_69 <= bright_gauss_ds_2_update_0_stage_68;
      bright_gauss_ds_2_update_0_stage_70 <= bright_gauss_ds_2_update_0_stage_69;
      bright_gauss_ds_2_update_0_stage_71 <= bright_gauss_ds_2_update_0_stage_70;
      bright_gauss_ds_2_update_0_stage_72 <= bright_gauss_ds_2_update_0_stage_71;
      bright_gauss_ds_2_update_0_stage_73 <= bright_gauss_ds_2_update_0_stage_72;
      bright_gauss_ds_2_update_0_stage_74 <= bright_gauss_ds_2_update_0_stage_73;
      bright_gauss_ds_2_update_0_stage_75 <= bright_gauss_ds_2_update_0_stage_74;
      bright_gauss_ds_2_update_0_stage_76 <= bright_gauss_ds_2_update_0_stage_75;
      bright_gauss_ds_2_update_0_stage_77 <= bright_gauss_ds_2_update_0_stage_76;
      bright_gauss_ds_2_update_0_stage_78 <= bright_gauss_ds_2_update_0_stage_77;
      bright_gauss_ds_2_update_0_stage_79 <= bright_gauss_ds_2_update_0_stage_78;
      bright_gauss_ds_2_update_0_stage_80 <= bright_gauss_ds_2_update_0_stage_79;
      bright_gauss_ds_2_update_0_stage_81 <= bright_gauss_ds_2_update_0_stage_80;
      bright_gauss_ds_2_update_0_stage_82 <= bright_gauss_ds_2_update_0_stage_81;
      bright_gauss_ds_2_update_0_stage_83 <= bright_gauss_ds_2_update_0_stage_82;
      bright_gauss_ds_2_update_0_stage_84 <= bright_gauss_ds_2_update_0_stage_83;
      bright_gauss_ds_2_update_0_stage_85 <= bright_gauss_ds_2_update_0_stage_84;
      bright_gauss_ds_2_update_0_stage_86 <= bright_gauss_ds_2_update_0_stage_85;
      bright_gauss_ds_2_update_0_stage_87 <= bright_gauss_ds_2_update_0_stage_86;
      bright_gauss_ds_2_update_0_stage_88 <= bright_gauss_ds_2_update_0_stage_87;
      bright_gauss_ds_2_update_0_stage_89 <= bright_gauss_ds_2_update_0_stage_88;
      bright_gauss_ds_2_update_0_stage_90 <= bright_gauss_ds_2_update_0_stage_89;
      bright_gauss_ds_2_update_0_stage_91 <= bright_gauss_ds_2_update_0_stage_90;
      bright_gauss_ds_2_update_0_stage_92 <= bright_gauss_ds_2_update_0_stage_91;
      bright_gauss_ds_2_update_0_stage_93 <= bright_gauss_ds_2_update_0_stage_92;
      bright_gauss_ds_2_update_0_stage_94 <= bright_gauss_ds_2_update_0_stage_93;
      bright_gauss_ds_2_update_0_stage_95 <= bright_gauss_ds_2_update_0_stage_94;
      bright_gauss_ds_2_update_0_stage_96 <= bright_gauss_ds_2_update_0_stage_95;
      bright_gauss_ds_2_update_0_stage_97 <= bright_gauss_ds_2_update_0_stage_96;
      bright_gauss_ds_2_update_0_stage_98 <= bright_gauss_ds_2_update_0_stage_97;
      bright_gauss_ds_2_update_0_stage_99 <= bright_gauss_ds_2_update_0_stage_98;
      bright_gauss_ds_2_update_0_stage_100 <= bright_gauss_ds_2_update_0_stage_99;
      bright_gauss_ds_2_update_0_stage_101 <= bright_gauss_ds_2_update_0_stage_100;
      bright_gauss_ds_2_update_0_stage_102 <= bright_gauss_ds_2_update_0_stage_101;
      bright_gauss_ds_2_update_0_stage_103 <= bright_gauss_ds_2_update_0_stage_102;
      bright_gauss_ds_2_update_0_stage_104 <= bright_gauss_ds_2_update_0_stage_103;
      bright_gauss_ds_2_update_0_stage_105 <= bright_gauss_ds_2_update_0_stage_104;
      bright_gauss_ds_2_update_0_stage_106 <= bright_gauss_ds_2_update_0_stage_105;
      bright_gauss_ds_2_update_0_stage_107 <= bright_gauss_ds_2_update_0_stage_106;
      bright_gauss_ds_2_update_0_stage_108 <= bright_gauss_ds_2_update_0_stage_107;
      bright_gauss_ds_2_update_0_stage_109 <= bright_gauss_ds_2_update_0_stage_108;
      bright_gauss_ds_2_update_0_stage_110 <= bright_gauss_ds_2_update_0_stage_109;
      bright_gauss_ds_2_update_0_stage_111 <= bright_gauss_ds_2_update_0_stage_110;
      bright_gauss_ds_2_update_0_stage_112 <= bright_gauss_ds_2_update_0_stage_111;
      bright_gauss_ds_2_update_0_stage_113 <= bright_gauss_ds_2_update_0_stage_112;
      bright_gauss_ds_2_update_0_stage_114 <= bright_gauss_ds_2_update_0_stage_113;
      bright_gauss_ds_2_update_0_stage_115 <= bright_gauss_ds_2_update_0_stage_114;
      bright_gauss_ds_2_update_0_stage_116 <= bright_gauss_ds_2_update_0_stage_115;
      bright_gauss_ds_2_update_0_stage_117 <= bright_gauss_ds_2_update_0_stage_116;
      bright_gauss_ds_2_update_0_stage_118 <= bright_gauss_ds_2_update_0_stage_117;
      bright_gauss_ds_2_update_0_stage_119 <= bright_gauss_ds_2_update_0_stage_118;
      bright_gauss_ds_2_update_0_stage_120 <= bright_gauss_ds_2_update_0_stage_119;
      bright_gauss_ds_2_update_0_stage_121 <= bright_gauss_ds_2_update_0_stage_120;
      bright_gauss_ds_2_update_0_stage_122 <= bright_gauss_ds_2_update_0_stage_121;
      bright_gauss_ds_2_update_0_stage_123 <= bright_gauss_ds_2_update_0_stage_122;
      bright_gauss_ds_2_update_0_stage_124 <= bright_gauss_ds_2_update_0_stage_123;
      bright_gauss_ds_2_update_0_stage_125 <= bright_gauss_ds_2_update_0_stage_124;
      bright_gauss_ds_2_update_0_stage_126 <= bright_gauss_ds_2_update_0_stage_125;
      bright_gauss_ds_2_update_0_stage_127 <= bright_gauss_ds_2_update_0_stage_126;
      bright_gauss_ds_2_update_0_stage_128 <= bright_gauss_ds_2_update_0_stage_127;
      bright_gauss_ds_2_update_0_stage_129 <= bright_gauss_ds_2_update_0_stage_128;
      bright_gauss_ds_2_update_0_stage_130 <= bright_gauss_ds_2_update_0_stage_129;
      bright_gauss_ds_2_update_0_stage_131 <= bright_gauss_ds_2_update_0_stage_130;
      bright_gauss_ds_2_update_0_stage_132 <= bright_gauss_ds_2_update_0_stage_131;
      bright_gauss_ds_2_update_0_stage_133 <= bright_gauss_ds_2_update_0_stage_132;
      bright_gauss_ds_2_update_0_stage_134 <= bright_gauss_ds_2_update_0_stage_133;
      bright_gauss_ds_2_update_0_stage_135 <= bright_gauss_ds_2_update_0_stage_134;
      bright_gauss_ds_2_update_0_stage_136 <= bright_gauss_ds_2_update_0_stage_135;
      bright_gauss_ds_2_update_0_stage_137 <= bright_gauss_ds_2_update_0_stage_136;
      bright_gauss_ds_2_update_0_stage_138 <= bright_gauss_ds_2_update_0_stage_137;
      bright_gauss_ds_2_update_0_stage_139 <= bright_gauss_ds_2_update_0_stage_138;
      bright_gauss_ds_2_update_0_stage_140 <= bright_gauss_ds_2_update_0_stage_139;
      bright_gauss_ds_2_update_0_stage_141 <= bright_gauss_ds_2_update_0_stage_140;
      bright_gauss_ds_2_update_0_stage_142 <= bright_gauss_ds_2_update_0_stage_141;
      bright_gauss_ds_2_update_0_stage_143 <= bright_gauss_ds_2_update_0_stage_142;
      bright_gauss_ds_2_update_0_stage_144 <= bright_gauss_ds_2_update_0_stage_143;
      bright_gauss_ds_2_update_0_stage_145 <= bright_gauss_ds_2_update_0_stage_144;
      bright_gauss_ds_2_update_0_stage_146 <= bright_gauss_ds_2_update_0_stage_145;
      bright_gauss_ds_2_update_0_stage_147 <= bright_gauss_ds_2_update_0_stage_146;
      bright_gauss_ds_2_update_0_stage_148 <= bright_gauss_ds_2_update_0_stage_147;
      bright_gauss_ds_2_update_0_stage_149 <= bright_gauss_ds_2_update_0_stage_148;
      bright_gauss_ds_2_update_0_stage_150 <= bright_gauss_ds_2_update_0_stage_149;
      bright_gauss_ds_2_update_0_stage_151 <= bright_gauss_ds_2_update_0_stage_150;
      bright_gauss_ds_2_update_0_stage_152 <= bright_gauss_ds_2_update_0_stage_151;
      bright_gauss_ds_2_update_0_stage_153 <= bright_gauss_ds_2_update_0_stage_152;
      bright_gauss_ds_2_update_0_stage_154 <= bright_gauss_ds_2_update_0_stage_153;
      bright_gauss_ds_2_update_0_stage_155 <= bright_gauss_ds_2_update_0_stage_154;
      bright_gauss_ds_2_update_0_stage_156 <= bright_gauss_ds_2_update_0_stage_155;
      bright_gauss_ds_2_update_0_stage_157 <= bright_gauss_ds_2_update_0_stage_156;
      bright_gauss_ds_2_update_0_stage_158 <= bright_gauss_ds_2_update_0_stage_157;
      bright_gauss_ds_2_update_0_stage_159 <= bright_gauss_ds_2_update_0_stage_158;
      bright_gauss_ds_2_update_0_stage_160 <= bright_gauss_ds_2_update_0_stage_159;
      bright_gauss_ds_2_update_0_stage_161 <= bright_gauss_ds_2_update_0_stage_160;
      bright_gauss_ds_2_update_0_stage_162 <= bright_gauss_ds_2_update_0_stage_161;
      bright_gauss_ds_2_update_0_stage_163 <= bright_gauss_ds_2_update_0_stage_162;
      bright_gauss_ds_2_update_0_stage_164 <= bright_gauss_ds_2_update_0_stage_163;
      bright_gauss_ds_2_update_0_stage_165 <= bright_gauss_ds_2_update_0_stage_164;
      bright_gauss_ds_2_update_0_stage_166 <= bright_gauss_ds_2_update_0_stage_165;
      bright_gauss_ds_2_update_0_stage_167 <= bright_gauss_ds_2_update_0_stage_166;
      bright_gauss_ds_2_update_0_stage_168 <= bright_gauss_ds_2_update_0_stage_167;
      bright_gauss_ds_2_update_0_stage_169 <= bright_gauss_ds_2_update_0_stage_168;
      bright_gauss_ds_2_update_0_stage_170 <= bright_gauss_ds_2_update_0_stage_169;
      bright_gauss_ds_2_update_0_stage_171 <= bright_gauss_ds_2_update_0_stage_170;
      bright_gauss_ds_2_update_0_stage_172 <= bright_gauss_ds_2_update_0_stage_171;
      bright_gauss_ds_2_update_0_stage_173 <= bright_gauss_ds_2_update_0_stage_172;
      bright_gauss_ds_2_update_0_stage_174 <= bright_gauss_ds_2_update_0_stage_173;
      bright_gauss_ds_2_update_0_stage_175 <= bright_gauss_ds_2_update_0_stage_174;
      bright_gauss_ds_2_update_0_stage_176 <= bright_gauss_ds_2_update_0_stage_175;
      bright_gauss_ds_2_update_0_stage_177 <= bright_gauss_ds_2_update_0_stage_176;
      bright_gauss_ds_2_update_0_stage_178 <= bright_gauss_ds_2_update_0_stage_177;
      bright_gauss_ds_2_update_0_stage_179 <= bright_gauss_ds_2_update_0_stage_178;
      bright_gauss_ds_2_update_0_stage_180 <= bright_gauss_ds_2_update_0_stage_179;
      bright_gauss_ds_2_update_0_stage_181 <= bright_gauss_ds_2_update_0_stage_180;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_58 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_59 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_58;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_60 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_59;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_61 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_60;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_62 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_61;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_63 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_62;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_64 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_63;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_65 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_64;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_66 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_65;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_67 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_66;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_68 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_67;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_69 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_68;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_70 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_69;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_71 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_70;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_72 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_71;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_73 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_72;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_74 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_73;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_75 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_74;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_76 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_75;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_77 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_76;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_78 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_77;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_79 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_78;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_80 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_79;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_81 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_80;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_82 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_81;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_83 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_82;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_84 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_83;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_85 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_84;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_86 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_85;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_87 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_86;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_88 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_87;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_89 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_88;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_90 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_89;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_91 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_90;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_92 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_91;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_93 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_92;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_94 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_93;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_95 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_94;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_96 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_95;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_97 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_96;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_98 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_97;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_99 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_98;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_100 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_99;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_101 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_100;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_102 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_101;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_103 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_102;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_104 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_103;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_105 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_104;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_106 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_105;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_107 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_106;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_108 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_107;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_109 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_108;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_110 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_109;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_111 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_110;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_112 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_111;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_113 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_112;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_114 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_113;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_115 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_114;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_116 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_115;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_117 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_116;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_118 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_117;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_119 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_118;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_120 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_119;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_121 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_120;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_122 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_121;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_123 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_122;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_124 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_123;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_125 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_124;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_126 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_125;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_127 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_126;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_128 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_127;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_129 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_128;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_130 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_129;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_131 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_130;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_132 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_131;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_133 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_132;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_134 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_133;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_135 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_134;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_136 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_135;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_137 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_136;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_138 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_137;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_139 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_138;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_140 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_139;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_141 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_140;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_142 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_141;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_143 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_142;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_144 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_143;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_145 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_144;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_146 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_145;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_147 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_146;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_148 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_147;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_149 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_148;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_150 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_149;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_151 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_150;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_152 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_151;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_153 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_152;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_154 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_153;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_155 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_154;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_156 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_155;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_157 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_156;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_158 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_157;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_159 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_158;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_160 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_159;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_161 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_160;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_162 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_161;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_163 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_162;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_164 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_163;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_165 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_164;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_166 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_165;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_167 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_166;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_168 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_167;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_169 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_168;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_170 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_169;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_171 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_170;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_172 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_171;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_173 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_172;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_174 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_173;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_175 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_174;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_176 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_175;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_177 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_176;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_178 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_177;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_179 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_178;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_180 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_179;
      bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_181 <= bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38_stage_180;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_51 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_52 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_51;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_53 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_52;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_54 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_53;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_55 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_54;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_56 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_55;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_57 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_56;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_58 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_57;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_59 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_58;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_60 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_59;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_61 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_60;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_62 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_61;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_63 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_62;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_64 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_63;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_65 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_64;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_66 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_65;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_67 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_66;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_68 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_67;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_69 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_68;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_70 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_69;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_71 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_70;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_72 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_71;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_73 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_72;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_74 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_73;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_75 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_74;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_76 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_75;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_77 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_76;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_78 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_77;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_79 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_78;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_80 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_79;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_81 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_80;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_82 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_81;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_83 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_82;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_84 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_83;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_85 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_84;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_86 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_85;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_87 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_86;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_88 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_87;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_89 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_88;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_90 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_89;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_91 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_90;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_92 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_91;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_93 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_92;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_94 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_93;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_95 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_94;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_96 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_95;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_97 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_96;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_98 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_97;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_99 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_98;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_100 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_99;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_101 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_100;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_102 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_101;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_103 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_102;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_104 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_103;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_105 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_104;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_106 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_105;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_107 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_106;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_108 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_107;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_109 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_108;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_110 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_109;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_111 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_110;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_112 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_111;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_113 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_112;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_114 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_113;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_115 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_114;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_116 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_115;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_117 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_116;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_118 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_117;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_119 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_118;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_120 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_119;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_121 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_120;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_122 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_121;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_123 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_122;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_124 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_123;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_125 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_124;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_126 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_125;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_127 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_126;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_128 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_127;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_129 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_128;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_130 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_129;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_131 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_130;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_132 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_131;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_133 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_132;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_134 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_133;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_135 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_134;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_136 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_135;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_137 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_136;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_138 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_137;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_139 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_138;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_140 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_139;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_141 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_140;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_142 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_141;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_143 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_142;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_144 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_143;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_145 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_144;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_146 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_145;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_147 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_146;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_148 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_147;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_149 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_148;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_150 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_149;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_151 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_150;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_152 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_151;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_153 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_152;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_154 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_153;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_155 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_154;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_156 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_155;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_157 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_156;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_158 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_157;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_159 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_158;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_160 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_159;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_161 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_160;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_162 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_161;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_163 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_162;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_164 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_163;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_165 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_164;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_166 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_165;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_167 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_166;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_168 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_167;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_169 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_168;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_170 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_169;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_171 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_170;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_172 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_171;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_173 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_172;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_174 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_173;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_175 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_174;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_176 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_175;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_177 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_176;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_178 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_177;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_179 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_178;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_180 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_179;
      bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_181 <= bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33_stage_180;
      bright_gauss_ds_3_update_0_stage_59 <= bright_gauss_ds_3_update_0;
      bright_gauss_ds_3_update_0_stage_60 <= bright_gauss_ds_3_update_0_stage_59;
      bright_gauss_ds_3_update_0_stage_61 <= bright_gauss_ds_3_update_0_stage_60;
      bright_gauss_ds_3_update_0_stage_62 <= bright_gauss_ds_3_update_0_stage_61;
      bright_gauss_ds_3_update_0_stage_63 <= bright_gauss_ds_3_update_0_stage_62;
      bright_gauss_ds_3_update_0_stage_64 <= bright_gauss_ds_3_update_0_stage_63;
      bright_gauss_ds_3_update_0_stage_65 <= bright_gauss_ds_3_update_0_stage_64;
      bright_gauss_ds_3_update_0_stage_66 <= bright_gauss_ds_3_update_0_stage_65;
      bright_gauss_ds_3_update_0_stage_67 <= bright_gauss_ds_3_update_0_stage_66;
      bright_gauss_ds_3_update_0_stage_68 <= bright_gauss_ds_3_update_0_stage_67;
      bright_gauss_ds_3_update_0_stage_69 <= bright_gauss_ds_3_update_0_stage_68;
      bright_gauss_ds_3_update_0_stage_70 <= bright_gauss_ds_3_update_0_stage_69;
      bright_gauss_ds_3_update_0_stage_71 <= bright_gauss_ds_3_update_0_stage_70;
      bright_gauss_ds_3_update_0_stage_72 <= bright_gauss_ds_3_update_0_stage_71;
      bright_gauss_ds_3_update_0_stage_73 <= bright_gauss_ds_3_update_0_stage_72;
      bright_gauss_ds_3_update_0_stage_74 <= bright_gauss_ds_3_update_0_stage_73;
      bright_gauss_ds_3_update_0_stage_75 <= bright_gauss_ds_3_update_0_stage_74;
      bright_gauss_ds_3_update_0_stage_76 <= bright_gauss_ds_3_update_0_stage_75;
      bright_gauss_ds_3_update_0_stage_77 <= bright_gauss_ds_3_update_0_stage_76;
      bright_gauss_ds_3_update_0_stage_78 <= bright_gauss_ds_3_update_0_stage_77;
      bright_gauss_ds_3_update_0_stage_79 <= bright_gauss_ds_3_update_0_stage_78;
      bright_gauss_ds_3_update_0_stage_80 <= bright_gauss_ds_3_update_0_stage_79;
      bright_gauss_ds_3_update_0_stage_81 <= bright_gauss_ds_3_update_0_stage_80;
      bright_gauss_ds_3_update_0_stage_82 <= bright_gauss_ds_3_update_0_stage_81;
      bright_gauss_ds_3_update_0_stage_83 <= bright_gauss_ds_3_update_0_stage_82;
      bright_gauss_ds_3_update_0_stage_84 <= bright_gauss_ds_3_update_0_stage_83;
      bright_gauss_ds_3_update_0_stage_85 <= bright_gauss_ds_3_update_0_stage_84;
      bright_gauss_ds_3_update_0_stage_86 <= bright_gauss_ds_3_update_0_stage_85;
      bright_gauss_ds_3_update_0_stage_87 <= bright_gauss_ds_3_update_0_stage_86;
      bright_gauss_ds_3_update_0_stage_88 <= bright_gauss_ds_3_update_0_stage_87;
      bright_gauss_ds_3_update_0_stage_89 <= bright_gauss_ds_3_update_0_stage_88;
      bright_gauss_ds_3_update_0_stage_90 <= bright_gauss_ds_3_update_0_stage_89;
      bright_gauss_ds_3_update_0_stage_91 <= bright_gauss_ds_3_update_0_stage_90;
      bright_gauss_ds_3_update_0_stage_92 <= bright_gauss_ds_3_update_0_stage_91;
      bright_gauss_ds_3_update_0_stage_93 <= bright_gauss_ds_3_update_0_stage_92;
      bright_gauss_ds_3_update_0_stage_94 <= bright_gauss_ds_3_update_0_stage_93;
      bright_gauss_ds_3_update_0_stage_95 <= bright_gauss_ds_3_update_0_stage_94;
      bright_gauss_ds_3_update_0_stage_96 <= bright_gauss_ds_3_update_0_stage_95;
      bright_gauss_ds_3_update_0_stage_97 <= bright_gauss_ds_3_update_0_stage_96;
      bright_gauss_ds_3_update_0_stage_98 <= bright_gauss_ds_3_update_0_stage_97;
      bright_gauss_ds_3_update_0_stage_99 <= bright_gauss_ds_3_update_0_stage_98;
      bright_gauss_ds_3_update_0_stage_100 <= bright_gauss_ds_3_update_0_stage_99;
      bright_gauss_ds_3_update_0_stage_101 <= bright_gauss_ds_3_update_0_stage_100;
      bright_gauss_ds_3_update_0_stage_102 <= bright_gauss_ds_3_update_0_stage_101;
      bright_gauss_ds_3_update_0_stage_103 <= bright_gauss_ds_3_update_0_stage_102;
      bright_gauss_ds_3_update_0_stage_104 <= bright_gauss_ds_3_update_0_stage_103;
      bright_gauss_ds_3_update_0_stage_105 <= bright_gauss_ds_3_update_0_stage_104;
      bright_gauss_ds_3_update_0_stage_106 <= bright_gauss_ds_3_update_0_stage_105;
      bright_gauss_ds_3_update_0_stage_107 <= bright_gauss_ds_3_update_0_stage_106;
      bright_gauss_ds_3_update_0_stage_108 <= bright_gauss_ds_3_update_0_stage_107;
      bright_gauss_ds_3_update_0_stage_109 <= bright_gauss_ds_3_update_0_stage_108;
      bright_gauss_ds_3_update_0_stage_110 <= bright_gauss_ds_3_update_0_stage_109;
      bright_gauss_ds_3_update_0_stage_111 <= bright_gauss_ds_3_update_0_stage_110;
      bright_gauss_ds_3_update_0_stage_112 <= bright_gauss_ds_3_update_0_stage_111;
      bright_gauss_ds_3_update_0_stage_113 <= bright_gauss_ds_3_update_0_stage_112;
      bright_gauss_ds_3_update_0_stage_114 <= bright_gauss_ds_3_update_0_stage_113;
      bright_gauss_ds_3_update_0_stage_115 <= bright_gauss_ds_3_update_0_stage_114;
      bright_gauss_ds_3_update_0_stage_116 <= bright_gauss_ds_3_update_0_stage_115;
      bright_gauss_ds_3_update_0_stage_117 <= bright_gauss_ds_3_update_0_stage_116;
      bright_gauss_ds_3_update_0_stage_118 <= bright_gauss_ds_3_update_0_stage_117;
      bright_gauss_ds_3_update_0_stage_119 <= bright_gauss_ds_3_update_0_stage_118;
      bright_gauss_ds_3_update_0_stage_120 <= bright_gauss_ds_3_update_0_stage_119;
      bright_gauss_ds_3_update_0_stage_121 <= bright_gauss_ds_3_update_0_stage_120;
      bright_gauss_ds_3_update_0_stage_122 <= bright_gauss_ds_3_update_0_stage_121;
      bright_gauss_ds_3_update_0_stage_123 <= bright_gauss_ds_3_update_0_stage_122;
      bright_gauss_ds_3_update_0_stage_124 <= bright_gauss_ds_3_update_0_stage_123;
      bright_gauss_ds_3_update_0_stage_125 <= bright_gauss_ds_3_update_0_stage_124;
      bright_gauss_ds_3_update_0_stage_126 <= bright_gauss_ds_3_update_0_stage_125;
      bright_gauss_ds_3_update_0_stage_127 <= bright_gauss_ds_3_update_0_stage_126;
      bright_gauss_ds_3_update_0_stage_128 <= bright_gauss_ds_3_update_0_stage_127;
      bright_gauss_ds_3_update_0_stage_129 <= bright_gauss_ds_3_update_0_stage_128;
      bright_gauss_ds_3_update_0_stage_130 <= bright_gauss_ds_3_update_0_stage_129;
      bright_gauss_ds_3_update_0_stage_131 <= bright_gauss_ds_3_update_0_stage_130;
      bright_gauss_ds_3_update_0_stage_132 <= bright_gauss_ds_3_update_0_stage_131;
      bright_gauss_ds_3_update_0_stage_133 <= bright_gauss_ds_3_update_0_stage_132;
      bright_gauss_ds_3_update_0_stage_134 <= bright_gauss_ds_3_update_0_stage_133;
      bright_gauss_ds_3_update_0_stage_135 <= bright_gauss_ds_3_update_0_stage_134;
      bright_gauss_ds_3_update_0_stage_136 <= bright_gauss_ds_3_update_0_stage_135;
      bright_gauss_ds_3_update_0_stage_137 <= bright_gauss_ds_3_update_0_stage_136;
      bright_gauss_ds_3_update_0_stage_138 <= bright_gauss_ds_3_update_0_stage_137;
      bright_gauss_ds_3_update_0_stage_139 <= bright_gauss_ds_3_update_0_stage_138;
      bright_gauss_ds_3_update_0_stage_140 <= bright_gauss_ds_3_update_0_stage_139;
      bright_gauss_ds_3_update_0_stage_141 <= bright_gauss_ds_3_update_0_stage_140;
      bright_gauss_ds_3_update_0_stage_142 <= bright_gauss_ds_3_update_0_stage_141;
      bright_gauss_ds_3_update_0_stage_143 <= bright_gauss_ds_3_update_0_stage_142;
      bright_gauss_ds_3_update_0_stage_144 <= bright_gauss_ds_3_update_0_stage_143;
      bright_gauss_ds_3_update_0_stage_145 <= bright_gauss_ds_3_update_0_stage_144;
      bright_gauss_ds_3_update_0_stage_146 <= bright_gauss_ds_3_update_0_stage_145;
      bright_gauss_ds_3_update_0_stage_147 <= bright_gauss_ds_3_update_0_stage_146;
      bright_gauss_ds_3_update_0_stage_148 <= bright_gauss_ds_3_update_0_stage_147;
      bright_gauss_ds_3_update_0_stage_149 <= bright_gauss_ds_3_update_0_stage_148;
      bright_gauss_ds_3_update_0_stage_150 <= bright_gauss_ds_3_update_0_stage_149;
      bright_gauss_ds_3_update_0_stage_151 <= bright_gauss_ds_3_update_0_stage_150;
      bright_gauss_ds_3_update_0_stage_152 <= bright_gauss_ds_3_update_0_stage_151;
      bright_gauss_ds_3_update_0_stage_153 <= bright_gauss_ds_3_update_0_stage_152;
      bright_gauss_ds_3_update_0_stage_154 <= bright_gauss_ds_3_update_0_stage_153;
      bright_gauss_ds_3_update_0_stage_155 <= bright_gauss_ds_3_update_0_stage_154;
      bright_gauss_ds_3_update_0_stage_156 <= bright_gauss_ds_3_update_0_stage_155;
      bright_gauss_ds_3_update_0_stage_157 <= bright_gauss_ds_3_update_0_stage_156;
      bright_gauss_ds_3_update_0_stage_158 <= bright_gauss_ds_3_update_0_stage_157;
      bright_gauss_ds_3_update_0_stage_159 <= bright_gauss_ds_3_update_0_stage_158;
      bright_gauss_ds_3_update_0_stage_160 <= bright_gauss_ds_3_update_0_stage_159;
      bright_gauss_ds_3_update_0_stage_161 <= bright_gauss_ds_3_update_0_stage_160;
      bright_gauss_ds_3_update_0_stage_162 <= bright_gauss_ds_3_update_0_stage_161;
      bright_gauss_ds_3_update_0_stage_163 <= bright_gauss_ds_3_update_0_stage_162;
      bright_gauss_ds_3_update_0_stage_164 <= bright_gauss_ds_3_update_0_stage_163;
      bright_gauss_ds_3_update_0_stage_165 <= bright_gauss_ds_3_update_0_stage_164;
      bright_gauss_ds_3_update_0_stage_166 <= bright_gauss_ds_3_update_0_stage_165;
      bright_gauss_ds_3_update_0_stage_167 <= bright_gauss_ds_3_update_0_stage_166;
      bright_gauss_ds_3_update_0_stage_168 <= bright_gauss_ds_3_update_0_stage_167;
      bright_gauss_ds_3_update_0_stage_169 <= bright_gauss_ds_3_update_0_stage_168;
      bright_gauss_ds_3_update_0_stage_170 <= bright_gauss_ds_3_update_0_stage_169;
      bright_gauss_ds_3_update_0_stage_171 <= bright_gauss_ds_3_update_0_stage_170;
      bright_gauss_ds_3_update_0_stage_172 <= bright_gauss_ds_3_update_0_stage_171;
      bright_gauss_ds_3_update_0_stage_173 <= bright_gauss_ds_3_update_0_stage_172;
      bright_gauss_ds_3_update_0_stage_174 <= bright_gauss_ds_3_update_0_stage_173;
      bright_gauss_ds_3_update_0_stage_175 <= bright_gauss_ds_3_update_0_stage_174;
      bright_gauss_ds_3_update_0_stage_176 <= bright_gauss_ds_3_update_0_stage_175;
      bright_gauss_ds_3_update_0_stage_177 <= bright_gauss_ds_3_update_0_stage_176;
      bright_gauss_ds_3_update_0_stage_178 <= bright_gauss_ds_3_update_0_stage_177;
      bright_gauss_ds_3_update_0_stage_179 <= bright_gauss_ds_3_update_0_stage_178;
      bright_gauss_ds_3_update_0_stage_180 <= bright_gauss_ds_3_update_0_stage_179;
      bright_gauss_ds_3_update_0_stage_181 <= bright_gauss_ds_3_update_0_stage_180;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_64 <= bright_bright_laplace_diff_0_update_0_read_read_42;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_65 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_64;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_66 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_65;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_67 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_66;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_68 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_67;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_69 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_68;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_70 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_69;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_71 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_70;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_72 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_71;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_73 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_72;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_74 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_73;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_75 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_74;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_76 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_75;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_77 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_76;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_78 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_77;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_79 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_78;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_80 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_79;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_81 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_80;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_82 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_81;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_83 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_82;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_84 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_83;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_85 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_84;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_86 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_85;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_87 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_86;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_88 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_87;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_89 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_88;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_90 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_89;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_91 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_90;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_92 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_91;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_93 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_92;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_94 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_93;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_95 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_94;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_96 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_95;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_97 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_96;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_98 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_97;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_99 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_98;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_100 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_99;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_101 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_100;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_102 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_101;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_103 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_102;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_104 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_103;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_105 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_104;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_106 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_105;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_107 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_106;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_108 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_107;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_109 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_108;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_110 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_109;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_111 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_110;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_112 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_111;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_113 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_112;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_114 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_113;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_115 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_114;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_116 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_115;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_117 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_116;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_118 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_117;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_119 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_118;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_120 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_119;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_121 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_120;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_122 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_121;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_123 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_122;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_124 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_123;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_125 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_124;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_126 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_125;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_127 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_126;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_128 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_127;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_129 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_128;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_130 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_129;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_131 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_130;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_132 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_131;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_133 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_132;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_134 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_133;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_135 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_134;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_136 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_135;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_137 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_136;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_138 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_137;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_139 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_138;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_140 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_139;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_141 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_140;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_142 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_141;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_143 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_142;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_144 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_143;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_145 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_144;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_146 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_145;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_147 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_146;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_148 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_147;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_149 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_148;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_150 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_149;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_151 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_150;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_152 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_151;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_153 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_152;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_154 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_153;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_155 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_154;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_156 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_155;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_157 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_156;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_158 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_157;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_159 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_158;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_160 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_159;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_161 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_160;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_162 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_161;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_163 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_162;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_164 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_163;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_165 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_164;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_166 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_165;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_167 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_166;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_168 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_167;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_169 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_168;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_170 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_169;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_171 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_170;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_172 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_171;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_173 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_172;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_174 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_173;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_175 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_174;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_176 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_175;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_177 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_176;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_178 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_177;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_179 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_178;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_180 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_179;
      bright_bright_laplace_diff_0_update_0_read_read_42_stage_181 <= bright_bright_laplace_diff_0_update_0_read_read_42_stage_180;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_65 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_66 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_65;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_67 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_66;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_68 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_67;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_69 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_68;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_70 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_69;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_71 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_70;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_72 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_71;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_73 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_72;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_74 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_73;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_75 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_74;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_76 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_75;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_77 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_76;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_78 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_77;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_79 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_78;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_80 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_79;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_81 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_80;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_82 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_81;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_83 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_82;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_84 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_83;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_85 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_84;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_86 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_85;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_87 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_86;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_88 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_87;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_89 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_88;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_90 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_89;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_91 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_90;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_92 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_91;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_93 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_92;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_94 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_93;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_95 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_94;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_96 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_95;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_97 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_96;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_98 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_97;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_99 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_98;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_100 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_99;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_101 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_100;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_102 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_101;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_103 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_102;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_104 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_103;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_105 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_104;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_106 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_105;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_107 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_106;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_108 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_107;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_109 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_108;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_110 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_109;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_111 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_110;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_112 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_111;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_113 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_112;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_114 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_113;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_115 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_114;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_116 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_115;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_117 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_116;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_118 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_117;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_119 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_118;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_120 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_119;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_121 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_120;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_122 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_121;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_123 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_122;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_124 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_123;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_125 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_124;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_126 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_125;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_127 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_126;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_128 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_127;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_129 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_128;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_130 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_129;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_131 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_130;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_132 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_131;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_133 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_132;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_134 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_133;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_135 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_134;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_136 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_135;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_137 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_136;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_138 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_137;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_139 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_138;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_140 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_139;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_141 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_140;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_142 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_141;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_143 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_142;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_144 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_143;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_145 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_144;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_146 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_145;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_147 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_146;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_148 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_147;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_149 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_148;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_150 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_149;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_151 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_150;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_152 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_151;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_153 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_152;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_154 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_153;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_155 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_154;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_156 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_155;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_157 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_156;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_158 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_157;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_159 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_158;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_160 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_159;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_161 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_160;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_162 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_161;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_163 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_162;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_164 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_163;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_165 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_164;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_166 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_165;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_167 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_166;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_168 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_167;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_169 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_168;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_170 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_169;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_171 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_170;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_172 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_171;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_173 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_172;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_174 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_173;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_175 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_174;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_176 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_175;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_177 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_176;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_178 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_177;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_179 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_178;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_180 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_179;
      bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_181 <= bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43_stage_180;
      bright_laplace_diff_0_update_0_stage_66 <= bright_laplace_diff_0_update_0;
      bright_laplace_diff_0_update_0_stage_67 <= bright_laplace_diff_0_update_0_stage_66;
      bright_laplace_diff_0_update_0_stage_68 <= bright_laplace_diff_0_update_0_stage_67;
      bright_laplace_diff_0_update_0_stage_69 <= bright_laplace_diff_0_update_0_stage_68;
      bright_laplace_diff_0_update_0_stage_70 <= bright_laplace_diff_0_update_0_stage_69;
      bright_laplace_diff_0_update_0_stage_71 <= bright_laplace_diff_0_update_0_stage_70;
      bright_laplace_diff_0_update_0_stage_72 <= bright_laplace_diff_0_update_0_stage_71;
      bright_laplace_diff_0_update_0_stage_73 <= bright_laplace_diff_0_update_0_stage_72;
      bright_laplace_diff_0_update_0_stage_74 <= bright_laplace_diff_0_update_0_stage_73;
      bright_laplace_diff_0_update_0_stage_75 <= bright_laplace_diff_0_update_0_stage_74;
      bright_laplace_diff_0_update_0_stage_76 <= bright_laplace_diff_0_update_0_stage_75;
      bright_laplace_diff_0_update_0_stage_77 <= bright_laplace_diff_0_update_0_stage_76;
      bright_laplace_diff_0_update_0_stage_78 <= bright_laplace_diff_0_update_0_stage_77;
      bright_laplace_diff_0_update_0_stage_79 <= bright_laplace_diff_0_update_0_stage_78;
      bright_laplace_diff_0_update_0_stage_80 <= bright_laplace_diff_0_update_0_stage_79;
      bright_laplace_diff_0_update_0_stage_81 <= bright_laplace_diff_0_update_0_stage_80;
      bright_laplace_diff_0_update_0_stage_82 <= bright_laplace_diff_0_update_0_stage_81;
      bright_laplace_diff_0_update_0_stage_83 <= bright_laplace_diff_0_update_0_stage_82;
      bright_laplace_diff_0_update_0_stage_84 <= bright_laplace_diff_0_update_0_stage_83;
      bright_laplace_diff_0_update_0_stage_85 <= bright_laplace_diff_0_update_0_stage_84;
      bright_laplace_diff_0_update_0_stage_86 <= bright_laplace_diff_0_update_0_stage_85;
      bright_laplace_diff_0_update_0_stage_87 <= bright_laplace_diff_0_update_0_stage_86;
      bright_laplace_diff_0_update_0_stage_88 <= bright_laplace_diff_0_update_0_stage_87;
      bright_laplace_diff_0_update_0_stage_89 <= bright_laplace_diff_0_update_0_stage_88;
      bright_laplace_diff_0_update_0_stage_90 <= bright_laplace_diff_0_update_0_stage_89;
      bright_laplace_diff_0_update_0_stage_91 <= bright_laplace_diff_0_update_0_stage_90;
      bright_laplace_diff_0_update_0_stage_92 <= bright_laplace_diff_0_update_0_stage_91;
      bright_laplace_diff_0_update_0_stage_93 <= bright_laplace_diff_0_update_0_stage_92;
      bright_laplace_diff_0_update_0_stage_94 <= bright_laplace_diff_0_update_0_stage_93;
      bright_laplace_diff_0_update_0_stage_95 <= bright_laplace_diff_0_update_0_stage_94;
      bright_laplace_diff_0_update_0_stage_96 <= bright_laplace_diff_0_update_0_stage_95;
      bright_laplace_diff_0_update_0_stage_97 <= bright_laplace_diff_0_update_0_stage_96;
      bright_laplace_diff_0_update_0_stage_98 <= bright_laplace_diff_0_update_0_stage_97;
      bright_laplace_diff_0_update_0_stage_99 <= bright_laplace_diff_0_update_0_stage_98;
      bright_laplace_diff_0_update_0_stage_100 <= bright_laplace_diff_0_update_0_stage_99;
      bright_laplace_diff_0_update_0_stage_101 <= bright_laplace_diff_0_update_0_stage_100;
      bright_laplace_diff_0_update_0_stage_102 <= bright_laplace_diff_0_update_0_stage_101;
      bright_laplace_diff_0_update_0_stage_103 <= bright_laplace_diff_0_update_0_stage_102;
      bright_laplace_diff_0_update_0_stage_104 <= bright_laplace_diff_0_update_0_stage_103;
      bright_laplace_diff_0_update_0_stage_105 <= bright_laplace_diff_0_update_0_stage_104;
      bright_laplace_diff_0_update_0_stage_106 <= bright_laplace_diff_0_update_0_stage_105;
      bright_laplace_diff_0_update_0_stage_107 <= bright_laplace_diff_0_update_0_stage_106;
      bright_laplace_diff_0_update_0_stage_108 <= bright_laplace_diff_0_update_0_stage_107;
      bright_laplace_diff_0_update_0_stage_109 <= bright_laplace_diff_0_update_0_stage_108;
      bright_laplace_diff_0_update_0_stage_110 <= bright_laplace_diff_0_update_0_stage_109;
      bright_laplace_diff_0_update_0_stage_111 <= bright_laplace_diff_0_update_0_stage_110;
      bright_laplace_diff_0_update_0_stage_112 <= bright_laplace_diff_0_update_0_stage_111;
      bright_laplace_diff_0_update_0_stage_113 <= bright_laplace_diff_0_update_0_stage_112;
      bright_laplace_diff_0_update_0_stage_114 <= bright_laplace_diff_0_update_0_stage_113;
      bright_laplace_diff_0_update_0_stage_115 <= bright_laplace_diff_0_update_0_stage_114;
      bright_laplace_diff_0_update_0_stage_116 <= bright_laplace_diff_0_update_0_stage_115;
      bright_laplace_diff_0_update_0_stage_117 <= bright_laplace_diff_0_update_0_stage_116;
      bright_laplace_diff_0_update_0_stage_118 <= bright_laplace_diff_0_update_0_stage_117;
      bright_laplace_diff_0_update_0_stage_119 <= bright_laplace_diff_0_update_0_stage_118;
      bright_laplace_diff_0_update_0_stage_120 <= bright_laplace_diff_0_update_0_stage_119;
      bright_laplace_diff_0_update_0_stage_121 <= bright_laplace_diff_0_update_0_stage_120;
      bright_laplace_diff_0_update_0_stage_122 <= bright_laplace_diff_0_update_0_stage_121;
      bright_laplace_diff_0_update_0_stage_123 <= bright_laplace_diff_0_update_0_stage_122;
      bright_laplace_diff_0_update_0_stage_124 <= bright_laplace_diff_0_update_0_stage_123;
      bright_laplace_diff_0_update_0_stage_125 <= bright_laplace_diff_0_update_0_stage_124;
      bright_laplace_diff_0_update_0_stage_126 <= bright_laplace_diff_0_update_0_stage_125;
      bright_laplace_diff_0_update_0_stage_127 <= bright_laplace_diff_0_update_0_stage_126;
      bright_laplace_diff_0_update_0_stage_128 <= bright_laplace_diff_0_update_0_stage_127;
      bright_laplace_diff_0_update_0_stage_129 <= bright_laplace_diff_0_update_0_stage_128;
      bright_laplace_diff_0_update_0_stage_130 <= bright_laplace_diff_0_update_0_stage_129;
      bright_laplace_diff_0_update_0_stage_131 <= bright_laplace_diff_0_update_0_stage_130;
      bright_laplace_diff_0_update_0_stage_132 <= bright_laplace_diff_0_update_0_stage_131;
      bright_laplace_diff_0_update_0_stage_133 <= bright_laplace_diff_0_update_0_stage_132;
      bright_laplace_diff_0_update_0_stage_134 <= bright_laplace_diff_0_update_0_stage_133;
      bright_laplace_diff_0_update_0_stage_135 <= bright_laplace_diff_0_update_0_stage_134;
      bright_laplace_diff_0_update_0_stage_136 <= bright_laplace_diff_0_update_0_stage_135;
      bright_laplace_diff_0_update_0_stage_137 <= bright_laplace_diff_0_update_0_stage_136;
      bright_laplace_diff_0_update_0_stage_138 <= bright_laplace_diff_0_update_0_stage_137;
      bright_laplace_diff_0_update_0_stage_139 <= bright_laplace_diff_0_update_0_stage_138;
      bright_laplace_diff_0_update_0_stage_140 <= bright_laplace_diff_0_update_0_stage_139;
      bright_laplace_diff_0_update_0_stage_141 <= bright_laplace_diff_0_update_0_stage_140;
      bright_laplace_diff_0_update_0_stage_142 <= bright_laplace_diff_0_update_0_stage_141;
      bright_laplace_diff_0_update_0_stage_143 <= bright_laplace_diff_0_update_0_stage_142;
      bright_laplace_diff_0_update_0_stage_144 <= bright_laplace_diff_0_update_0_stage_143;
      bright_laplace_diff_0_update_0_stage_145 <= bright_laplace_diff_0_update_0_stage_144;
      bright_laplace_diff_0_update_0_stage_146 <= bright_laplace_diff_0_update_0_stage_145;
      bright_laplace_diff_0_update_0_stage_147 <= bright_laplace_diff_0_update_0_stage_146;
      bright_laplace_diff_0_update_0_stage_148 <= bright_laplace_diff_0_update_0_stage_147;
      bright_laplace_diff_0_update_0_stage_149 <= bright_laplace_diff_0_update_0_stage_148;
      bright_laplace_diff_0_update_0_stage_150 <= bright_laplace_diff_0_update_0_stage_149;
      bright_laplace_diff_0_update_0_stage_151 <= bright_laplace_diff_0_update_0_stage_150;
      bright_laplace_diff_0_update_0_stage_152 <= bright_laplace_diff_0_update_0_stage_151;
      bright_laplace_diff_0_update_0_stage_153 <= bright_laplace_diff_0_update_0_stage_152;
      bright_laplace_diff_0_update_0_stage_154 <= bright_laplace_diff_0_update_0_stage_153;
      bright_laplace_diff_0_update_0_stage_155 <= bright_laplace_diff_0_update_0_stage_154;
      bright_laplace_diff_0_update_0_stage_156 <= bright_laplace_diff_0_update_0_stage_155;
      bright_laplace_diff_0_update_0_stage_157 <= bright_laplace_diff_0_update_0_stage_156;
      bright_laplace_diff_0_update_0_stage_158 <= bright_laplace_diff_0_update_0_stage_157;
      bright_laplace_diff_0_update_0_stage_159 <= bright_laplace_diff_0_update_0_stage_158;
      bright_laplace_diff_0_update_0_stage_160 <= bright_laplace_diff_0_update_0_stage_159;
      bright_laplace_diff_0_update_0_stage_161 <= bright_laplace_diff_0_update_0_stage_160;
      bright_laplace_diff_0_update_0_stage_162 <= bright_laplace_diff_0_update_0_stage_161;
      bright_laplace_diff_0_update_0_stage_163 <= bright_laplace_diff_0_update_0_stage_162;
      bright_laplace_diff_0_update_0_stage_164 <= bright_laplace_diff_0_update_0_stage_163;
      bright_laplace_diff_0_update_0_stage_165 <= bright_laplace_diff_0_update_0_stage_164;
      bright_laplace_diff_0_update_0_stage_166 <= bright_laplace_diff_0_update_0_stage_165;
      bright_laplace_diff_0_update_0_stage_167 <= bright_laplace_diff_0_update_0_stage_166;
      bright_laplace_diff_0_update_0_stage_168 <= bright_laplace_diff_0_update_0_stage_167;
      bright_laplace_diff_0_update_0_stage_169 <= bright_laplace_diff_0_update_0_stage_168;
      bright_laplace_diff_0_update_0_stage_170 <= bright_laplace_diff_0_update_0_stage_169;
      bright_laplace_diff_0_update_0_stage_171 <= bright_laplace_diff_0_update_0_stage_170;
      bright_laplace_diff_0_update_0_stage_172 <= bright_laplace_diff_0_update_0_stage_171;
      bright_laplace_diff_0_update_0_stage_173 <= bright_laplace_diff_0_update_0_stage_172;
      bright_laplace_diff_0_update_0_stage_174 <= bright_laplace_diff_0_update_0_stage_173;
      bright_laplace_diff_0_update_0_stage_175 <= bright_laplace_diff_0_update_0_stage_174;
      bright_laplace_diff_0_update_0_stage_176 <= bright_laplace_diff_0_update_0_stage_175;
      bright_laplace_diff_0_update_0_stage_177 <= bright_laplace_diff_0_update_0_stage_176;
      bright_laplace_diff_0_update_0_stage_178 <= bright_laplace_diff_0_update_0_stage_177;
      bright_laplace_diff_0_update_0_stage_179 <= bright_laplace_diff_0_update_0_stage_178;
      bright_laplace_diff_0_update_0_stage_180 <= bright_laplace_diff_0_update_0_stage_179;
      bright_laplace_diff_0_update_0_stage_181 <= bright_laplace_diff_0_update_0_stage_180;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_67 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_68 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_67;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_69 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_68;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_70 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_69;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_71 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_70;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_72 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_71;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_73 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_72;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_74 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_73;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_75 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_74;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_76 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_75;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_77 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_76;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_78 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_77;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_79 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_78;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_80 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_79;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_81 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_80;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_82 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_81;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_83 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_82;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_84 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_83;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_85 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_84;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_86 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_85;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_87 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_86;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_88 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_87;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_89 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_88;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_90 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_89;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_91 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_90;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_92 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_91;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_93 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_92;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_94 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_93;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_95 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_94;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_96 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_95;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_97 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_96;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_98 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_97;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_99 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_98;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_100 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_99;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_101 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_100;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_102 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_101;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_103 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_102;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_104 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_103;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_105 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_104;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_106 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_105;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_107 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_106;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_108 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_107;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_109 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_108;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_110 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_109;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_111 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_110;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_112 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_111;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_113 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_112;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_114 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_113;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_115 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_114;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_116 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_115;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_117 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_116;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_118 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_117;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_119 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_118;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_120 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_119;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_121 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_120;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_122 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_121;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_123 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_122;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_124 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_123;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_125 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_124;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_126 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_125;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_127 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_126;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_128 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_127;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_129 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_128;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_130 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_129;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_131 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_130;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_132 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_131;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_133 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_132;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_134 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_133;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_135 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_134;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_136 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_135;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_137 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_136;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_138 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_137;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_139 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_138;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_140 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_139;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_141 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_140;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_142 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_141;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_143 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_142;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_144 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_143;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_145 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_144;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_146 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_145;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_147 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_146;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_148 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_147;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_149 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_148;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_150 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_149;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_151 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_150;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_152 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_151;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_153 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_152;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_154 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_153;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_155 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_154;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_156 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_155;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_157 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_156;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_158 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_157;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_159 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_158;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_160 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_159;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_161 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_160;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_162 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_161;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_163 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_162;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_164 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_163;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_165 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_164;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_166 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_165;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_167 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_166;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_168 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_167;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_169 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_168;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_170 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_169;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_171 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_170;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_172 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_171;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_173 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_172;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_174 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_173;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_175 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_174;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_176 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_175;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_177 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_176;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_178 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_177;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_179 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_178;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_180 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_179;
      bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_181 <= bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44_stage_180;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_72 <= bright_weights_bright_weights_normed_update_0_read_read_48;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_73 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_72;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_74 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_73;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_75 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_74;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_76 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_75;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_77 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_76;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_78 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_77;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_79 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_78;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_80 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_79;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_81 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_80;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_82 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_81;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_83 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_82;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_84 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_83;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_85 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_84;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_86 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_85;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_87 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_86;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_88 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_87;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_89 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_88;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_90 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_89;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_91 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_90;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_92 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_91;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_93 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_92;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_94 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_93;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_95 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_94;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_96 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_95;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_97 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_96;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_98 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_97;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_99 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_98;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_100 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_99;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_101 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_100;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_102 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_101;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_103 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_102;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_104 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_103;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_105 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_104;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_106 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_105;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_107 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_106;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_108 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_107;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_109 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_108;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_110 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_109;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_111 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_110;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_112 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_111;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_113 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_112;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_114 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_113;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_115 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_114;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_116 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_115;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_117 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_116;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_118 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_117;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_119 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_118;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_120 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_119;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_121 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_120;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_122 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_121;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_123 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_122;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_124 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_123;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_125 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_124;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_126 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_125;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_127 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_126;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_128 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_127;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_129 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_128;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_130 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_129;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_131 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_130;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_132 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_131;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_133 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_132;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_134 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_133;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_135 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_134;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_136 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_135;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_137 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_136;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_138 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_137;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_139 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_138;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_140 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_139;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_141 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_140;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_142 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_141;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_143 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_142;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_144 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_143;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_145 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_144;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_146 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_145;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_147 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_146;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_148 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_147;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_149 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_148;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_150 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_149;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_151 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_150;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_152 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_151;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_153 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_152;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_154 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_153;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_155 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_154;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_156 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_155;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_157 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_156;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_158 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_157;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_159 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_158;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_160 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_159;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_161 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_160;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_162 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_161;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_163 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_162;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_164 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_163;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_165 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_164;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_166 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_165;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_167 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_166;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_168 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_167;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_169 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_168;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_170 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_169;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_171 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_170;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_172 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_171;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_173 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_172;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_174 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_173;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_175 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_174;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_176 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_175;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_177 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_176;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_178 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_177;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_179 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_178;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_180 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_179;
      bright_weights_bright_weights_normed_update_0_read_read_48_stage_181 <= bright_weights_bright_weights_normed_update_0_read_read_48_stage_180;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_73 <= weight_sums_bright_weights_normed_update_0_read_read_49;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_74 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_73;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_75 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_74;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_76 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_75;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_77 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_76;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_78 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_77;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_79 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_78;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_80 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_79;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_81 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_80;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_82 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_81;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_83 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_82;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_84 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_83;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_85 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_84;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_86 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_85;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_87 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_86;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_88 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_87;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_89 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_88;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_90 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_89;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_91 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_90;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_92 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_91;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_93 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_92;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_94 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_93;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_95 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_94;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_96 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_95;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_97 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_96;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_98 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_97;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_99 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_98;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_100 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_99;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_101 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_100;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_102 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_101;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_103 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_102;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_104 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_103;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_105 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_104;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_106 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_105;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_107 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_106;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_108 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_107;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_109 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_108;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_110 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_109;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_111 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_110;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_112 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_111;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_113 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_112;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_114 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_113;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_115 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_114;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_116 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_115;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_117 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_116;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_118 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_117;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_119 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_118;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_120 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_119;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_121 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_120;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_122 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_121;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_123 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_122;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_124 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_123;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_125 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_124;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_126 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_125;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_127 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_126;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_128 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_127;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_129 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_128;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_130 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_129;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_131 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_130;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_132 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_131;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_133 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_132;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_134 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_133;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_135 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_134;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_136 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_135;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_137 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_136;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_138 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_137;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_139 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_138;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_140 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_139;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_141 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_140;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_142 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_141;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_143 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_142;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_144 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_143;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_145 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_144;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_146 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_145;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_147 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_146;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_148 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_147;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_149 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_148;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_150 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_149;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_151 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_150;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_152 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_151;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_153 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_152;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_154 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_153;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_155 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_154;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_156 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_155;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_157 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_156;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_158 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_157;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_159 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_158;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_160 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_159;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_161 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_160;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_162 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_161;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_163 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_162;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_164 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_163;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_165 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_164;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_166 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_165;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_167 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_166;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_168 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_167;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_169 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_168;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_170 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_169;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_171 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_170;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_172 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_171;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_173 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_172;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_174 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_173;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_175 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_174;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_176 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_175;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_177 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_176;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_178 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_177;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_179 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_178;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_180 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_179;
      weight_sums_bright_weights_normed_update_0_read_read_49_stage_181 <= weight_sums_bright_weights_normed_update_0_read_read_49_stage_180;
      bright_weights_normed_update_0_stage_74 <= bright_weights_normed_update_0;
      bright_weights_normed_update_0_stage_75 <= bright_weights_normed_update_0_stage_74;
      bright_weights_normed_update_0_stage_76 <= bright_weights_normed_update_0_stage_75;
      bright_weights_normed_update_0_stage_77 <= bright_weights_normed_update_0_stage_76;
      bright_weights_normed_update_0_stage_78 <= bright_weights_normed_update_0_stage_77;
      bright_weights_normed_update_0_stage_79 <= bright_weights_normed_update_0_stage_78;
      bright_weights_normed_update_0_stage_80 <= bright_weights_normed_update_0_stage_79;
      bright_weights_normed_update_0_stage_81 <= bright_weights_normed_update_0_stage_80;
      bright_weights_normed_update_0_stage_82 <= bright_weights_normed_update_0_stage_81;
      bright_weights_normed_update_0_stage_83 <= bright_weights_normed_update_0_stage_82;
      bright_weights_normed_update_0_stage_84 <= bright_weights_normed_update_0_stage_83;
      bright_weights_normed_update_0_stage_85 <= bright_weights_normed_update_0_stage_84;
      bright_weights_normed_update_0_stage_86 <= bright_weights_normed_update_0_stage_85;
      bright_weights_normed_update_0_stage_87 <= bright_weights_normed_update_0_stage_86;
      bright_weights_normed_update_0_stage_88 <= bright_weights_normed_update_0_stage_87;
      bright_weights_normed_update_0_stage_89 <= bright_weights_normed_update_0_stage_88;
      bright_weights_normed_update_0_stage_90 <= bright_weights_normed_update_0_stage_89;
      bright_weights_normed_update_0_stage_91 <= bright_weights_normed_update_0_stage_90;
      bright_weights_normed_update_0_stage_92 <= bright_weights_normed_update_0_stage_91;
      bright_weights_normed_update_0_stage_93 <= bright_weights_normed_update_0_stage_92;
      bright_weights_normed_update_0_stage_94 <= bright_weights_normed_update_0_stage_93;
      bright_weights_normed_update_0_stage_95 <= bright_weights_normed_update_0_stage_94;
      bright_weights_normed_update_0_stage_96 <= bright_weights_normed_update_0_stage_95;
      bright_weights_normed_update_0_stage_97 <= bright_weights_normed_update_0_stage_96;
      bright_weights_normed_update_0_stage_98 <= bright_weights_normed_update_0_stage_97;
      bright_weights_normed_update_0_stage_99 <= bright_weights_normed_update_0_stage_98;
      bright_weights_normed_update_0_stage_100 <= bright_weights_normed_update_0_stage_99;
      bright_weights_normed_update_0_stage_101 <= bright_weights_normed_update_0_stage_100;
      bright_weights_normed_update_0_stage_102 <= bright_weights_normed_update_0_stage_101;
      bright_weights_normed_update_0_stage_103 <= bright_weights_normed_update_0_stage_102;
      bright_weights_normed_update_0_stage_104 <= bright_weights_normed_update_0_stage_103;
      bright_weights_normed_update_0_stage_105 <= bright_weights_normed_update_0_stage_104;
      bright_weights_normed_update_0_stage_106 <= bright_weights_normed_update_0_stage_105;
      bright_weights_normed_update_0_stage_107 <= bright_weights_normed_update_0_stage_106;
      bright_weights_normed_update_0_stage_108 <= bright_weights_normed_update_0_stage_107;
      bright_weights_normed_update_0_stage_109 <= bright_weights_normed_update_0_stage_108;
      bright_weights_normed_update_0_stage_110 <= bright_weights_normed_update_0_stage_109;
      bright_weights_normed_update_0_stage_111 <= bright_weights_normed_update_0_stage_110;
      bright_weights_normed_update_0_stage_112 <= bright_weights_normed_update_0_stage_111;
      bright_weights_normed_update_0_stage_113 <= bright_weights_normed_update_0_stage_112;
      bright_weights_normed_update_0_stage_114 <= bright_weights_normed_update_0_stage_113;
      bright_weights_normed_update_0_stage_115 <= bright_weights_normed_update_0_stage_114;
      bright_weights_normed_update_0_stage_116 <= bright_weights_normed_update_0_stage_115;
      bright_weights_normed_update_0_stage_117 <= bright_weights_normed_update_0_stage_116;
      bright_weights_normed_update_0_stage_118 <= bright_weights_normed_update_0_stage_117;
      bright_weights_normed_update_0_stage_119 <= bright_weights_normed_update_0_stage_118;
      bright_weights_normed_update_0_stage_120 <= bright_weights_normed_update_0_stage_119;
      bright_weights_normed_update_0_stage_121 <= bright_weights_normed_update_0_stage_120;
      bright_weights_normed_update_0_stage_122 <= bright_weights_normed_update_0_stage_121;
      bright_weights_normed_update_0_stage_123 <= bright_weights_normed_update_0_stage_122;
      bright_weights_normed_update_0_stage_124 <= bright_weights_normed_update_0_stage_123;
      bright_weights_normed_update_0_stage_125 <= bright_weights_normed_update_0_stage_124;
      bright_weights_normed_update_0_stage_126 <= bright_weights_normed_update_0_stage_125;
      bright_weights_normed_update_0_stage_127 <= bright_weights_normed_update_0_stage_126;
      bright_weights_normed_update_0_stage_128 <= bright_weights_normed_update_0_stage_127;
      bright_weights_normed_update_0_stage_129 <= bright_weights_normed_update_0_stage_128;
      bright_weights_normed_update_0_stage_130 <= bright_weights_normed_update_0_stage_129;
      bright_weights_normed_update_0_stage_131 <= bright_weights_normed_update_0_stage_130;
      bright_weights_normed_update_0_stage_132 <= bright_weights_normed_update_0_stage_131;
      bright_weights_normed_update_0_stage_133 <= bright_weights_normed_update_0_stage_132;
      bright_weights_normed_update_0_stage_134 <= bright_weights_normed_update_0_stage_133;
      bright_weights_normed_update_0_stage_135 <= bright_weights_normed_update_0_stage_134;
      bright_weights_normed_update_0_stage_136 <= bright_weights_normed_update_0_stage_135;
      bright_weights_normed_update_0_stage_137 <= bright_weights_normed_update_0_stage_136;
      bright_weights_normed_update_0_stage_138 <= bright_weights_normed_update_0_stage_137;
      bright_weights_normed_update_0_stage_139 <= bright_weights_normed_update_0_stage_138;
      bright_weights_normed_update_0_stage_140 <= bright_weights_normed_update_0_stage_139;
      bright_weights_normed_update_0_stage_141 <= bright_weights_normed_update_0_stage_140;
      bright_weights_normed_update_0_stage_142 <= bright_weights_normed_update_0_stage_141;
      bright_weights_normed_update_0_stage_143 <= bright_weights_normed_update_0_stage_142;
      bright_weights_normed_update_0_stage_144 <= bright_weights_normed_update_0_stage_143;
      bright_weights_normed_update_0_stage_145 <= bright_weights_normed_update_0_stage_144;
      bright_weights_normed_update_0_stage_146 <= bright_weights_normed_update_0_stage_145;
      bright_weights_normed_update_0_stage_147 <= bright_weights_normed_update_0_stage_146;
      bright_weights_normed_update_0_stage_148 <= bright_weights_normed_update_0_stage_147;
      bright_weights_normed_update_0_stage_149 <= bright_weights_normed_update_0_stage_148;
      bright_weights_normed_update_0_stage_150 <= bright_weights_normed_update_0_stage_149;
      bright_weights_normed_update_0_stage_151 <= bright_weights_normed_update_0_stage_150;
      bright_weights_normed_update_0_stage_152 <= bright_weights_normed_update_0_stage_151;
      bright_weights_normed_update_0_stage_153 <= bright_weights_normed_update_0_stage_152;
      bright_weights_normed_update_0_stage_154 <= bright_weights_normed_update_0_stage_153;
      bright_weights_normed_update_0_stage_155 <= bright_weights_normed_update_0_stage_154;
      bright_weights_normed_update_0_stage_156 <= bright_weights_normed_update_0_stage_155;
      bright_weights_normed_update_0_stage_157 <= bright_weights_normed_update_0_stage_156;
      bright_weights_normed_update_0_stage_158 <= bright_weights_normed_update_0_stage_157;
      bright_weights_normed_update_0_stage_159 <= bright_weights_normed_update_0_stage_158;
      bright_weights_normed_update_0_stage_160 <= bright_weights_normed_update_0_stage_159;
      bright_weights_normed_update_0_stage_161 <= bright_weights_normed_update_0_stage_160;
      bright_weights_normed_update_0_stage_162 <= bright_weights_normed_update_0_stage_161;
      bright_weights_normed_update_0_stage_163 <= bright_weights_normed_update_0_stage_162;
      bright_weights_normed_update_0_stage_164 <= bright_weights_normed_update_0_stage_163;
      bright_weights_normed_update_0_stage_165 <= bright_weights_normed_update_0_stage_164;
      bright_weights_normed_update_0_stage_166 <= bright_weights_normed_update_0_stage_165;
      bright_weights_normed_update_0_stage_167 <= bright_weights_normed_update_0_stage_166;
      bright_weights_normed_update_0_stage_168 <= bright_weights_normed_update_0_stage_167;
      bright_weights_normed_update_0_stage_169 <= bright_weights_normed_update_0_stage_168;
      bright_weights_normed_update_0_stage_170 <= bright_weights_normed_update_0_stage_169;
      bright_weights_normed_update_0_stage_171 <= bright_weights_normed_update_0_stage_170;
      bright_weights_normed_update_0_stage_172 <= bright_weights_normed_update_0_stage_171;
      bright_weights_normed_update_0_stage_173 <= bright_weights_normed_update_0_stage_172;
      bright_weights_normed_update_0_stage_174 <= bright_weights_normed_update_0_stage_173;
      bright_weights_normed_update_0_stage_175 <= bright_weights_normed_update_0_stage_174;
      bright_weights_normed_update_0_stage_176 <= bright_weights_normed_update_0_stage_175;
      bright_weights_normed_update_0_stage_177 <= bright_weights_normed_update_0_stage_176;
      bright_weights_normed_update_0_stage_178 <= bright_weights_normed_update_0_stage_177;
      bright_weights_normed_update_0_stage_179 <= bright_weights_normed_update_0_stage_178;
      bright_weights_normed_update_0_stage_180 <= bright_weights_normed_update_0_stage_179;
      bright_weights_normed_update_0_stage_181 <= bright_weights_normed_update_0_stage_180;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_75 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_76 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_75;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_77 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_76;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_78 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_77;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_79 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_78;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_80 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_79;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_81 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_80;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_82 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_81;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_83 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_82;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_84 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_83;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_85 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_84;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_86 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_85;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_87 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_86;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_88 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_87;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_89 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_88;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_90 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_89;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_91 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_90;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_92 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_91;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_93 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_92;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_94 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_93;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_95 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_94;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_96 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_95;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_97 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_96;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_98 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_97;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_99 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_98;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_100 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_99;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_101 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_100;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_102 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_101;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_103 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_102;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_104 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_103;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_105 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_104;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_106 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_105;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_107 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_106;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_108 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_107;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_109 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_108;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_110 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_109;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_111 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_110;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_112 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_111;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_113 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_112;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_114 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_113;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_115 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_114;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_116 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_115;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_117 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_116;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_118 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_117;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_119 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_118;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_120 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_119;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_121 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_120;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_122 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_121;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_123 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_122;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_124 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_123;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_125 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_124;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_126 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_125;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_127 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_126;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_128 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_127;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_129 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_128;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_130 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_129;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_131 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_130;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_132 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_131;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_133 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_132;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_134 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_133;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_135 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_134;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_136 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_135;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_137 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_136;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_138 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_137;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_139 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_138;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_140 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_139;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_141 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_140;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_142 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_141;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_143 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_142;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_144 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_143;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_145 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_144;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_146 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_145;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_147 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_146;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_148 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_147;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_149 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_148;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_150 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_149;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_151 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_150;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_152 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_151;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_153 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_152;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_154 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_153;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_155 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_154;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_156 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_155;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_157 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_156;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_158 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_157;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_159 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_158;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_160 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_159;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_161 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_160;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_162 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_161;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_163 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_162;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_164 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_163;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_165 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_164;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_166 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_165;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_167 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_166;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_168 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_167;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_169 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_168;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_170 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_169;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_171 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_170;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_172 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_171;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_173 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_172;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_174 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_173;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_175 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_174;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_176 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_175;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_177 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_176;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_178 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_177;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_179 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_178;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_180 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_179;
      bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_181 <= bright_weights_normed_bright_weights_normed_update_0_write_write_50_stage_180;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_79 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_80 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_79;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_81 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_80;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_82 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_81;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_83 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_82;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_84 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_83;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_85 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_84;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_86 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_85;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_87 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_86;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_88 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_87;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_89 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_88;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_90 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_89;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_91 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_90;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_92 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_91;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_93 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_92;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_94 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_93;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_95 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_94;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_96 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_95;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_97 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_96;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_98 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_97;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_99 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_98;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_100 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_99;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_101 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_100;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_102 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_101;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_103 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_102;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_104 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_103;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_105 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_104;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_106 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_105;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_107 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_106;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_108 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_107;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_109 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_108;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_110 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_109;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_111 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_110;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_112 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_111;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_113 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_112;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_114 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_113;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_115 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_114;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_116 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_115;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_117 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_116;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_118 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_117;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_119 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_118;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_120 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_119;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_121 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_120;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_122 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_121;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_123 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_122;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_124 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_123;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_125 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_124;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_126 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_125;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_127 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_126;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_128 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_127;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_129 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_128;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_130 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_129;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_131 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_130;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_132 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_131;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_133 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_132;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_134 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_133;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_135 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_134;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_136 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_135;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_137 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_136;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_138 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_137;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_139 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_138;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_140 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_139;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_141 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_140;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_142 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_141;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_143 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_142;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_144 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_143;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_145 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_144;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_146 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_145;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_147 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_146;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_148 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_147;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_149 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_148;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_150 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_149;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_151 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_150;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_152 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_151;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_153 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_152;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_154 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_153;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_155 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_154;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_156 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_155;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_157 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_156;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_158 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_157;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_159 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_158;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_160 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_159;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_161 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_160;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_162 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_161;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_163 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_162;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_164 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_163;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_165 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_164;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_166 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_165;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_167 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_166;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_168 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_167;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_169 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_168;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_170 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_169;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_171 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_170;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_172 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_171;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_173 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_172;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_174 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_173;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_175 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_174;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_176 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_175;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_177 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_176;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_178 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_177;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_179 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_178;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_180 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_179;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_181 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53_stage_180;
      dark_weights_normed_gauss_ds_1_update_0_stage_80 <= dark_weights_normed_gauss_ds_1_update_0;
      dark_weights_normed_gauss_ds_1_update_0_stage_81 <= dark_weights_normed_gauss_ds_1_update_0_stage_80;
      dark_weights_normed_gauss_ds_1_update_0_stage_82 <= dark_weights_normed_gauss_ds_1_update_0_stage_81;
      dark_weights_normed_gauss_ds_1_update_0_stage_83 <= dark_weights_normed_gauss_ds_1_update_0_stage_82;
      dark_weights_normed_gauss_ds_1_update_0_stage_84 <= dark_weights_normed_gauss_ds_1_update_0_stage_83;
      dark_weights_normed_gauss_ds_1_update_0_stage_85 <= dark_weights_normed_gauss_ds_1_update_0_stage_84;
      dark_weights_normed_gauss_ds_1_update_0_stage_86 <= dark_weights_normed_gauss_ds_1_update_0_stage_85;
      dark_weights_normed_gauss_ds_1_update_0_stage_87 <= dark_weights_normed_gauss_ds_1_update_0_stage_86;
      dark_weights_normed_gauss_ds_1_update_0_stage_88 <= dark_weights_normed_gauss_ds_1_update_0_stage_87;
      dark_weights_normed_gauss_ds_1_update_0_stage_89 <= dark_weights_normed_gauss_ds_1_update_0_stage_88;
      dark_weights_normed_gauss_ds_1_update_0_stage_90 <= dark_weights_normed_gauss_ds_1_update_0_stage_89;
      dark_weights_normed_gauss_ds_1_update_0_stage_91 <= dark_weights_normed_gauss_ds_1_update_0_stage_90;
      dark_weights_normed_gauss_ds_1_update_0_stage_92 <= dark_weights_normed_gauss_ds_1_update_0_stage_91;
      dark_weights_normed_gauss_ds_1_update_0_stage_93 <= dark_weights_normed_gauss_ds_1_update_0_stage_92;
      dark_weights_normed_gauss_ds_1_update_0_stage_94 <= dark_weights_normed_gauss_ds_1_update_0_stage_93;
      dark_weights_normed_gauss_ds_1_update_0_stage_95 <= dark_weights_normed_gauss_ds_1_update_0_stage_94;
      dark_weights_normed_gauss_ds_1_update_0_stage_96 <= dark_weights_normed_gauss_ds_1_update_0_stage_95;
      dark_weights_normed_gauss_ds_1_update_0_stage_97 <= dark_weights_normed_gauss_ds_1_update_0_stage_96;
      dark_weights_normed_gauss_ds_1_update_0_stage_98 <= dark_weights_normed_gauss_ds_1_update_0_stage_97;
      dark_weights_normed_gauss_ds_1_update_0_stage_99 <= dark_weights_normed_gauss_ds_1_update_0_stage_98;
      dark_weights_normed_gauss_ds_1_update_0_stage_100 <= dark_weights_normed_gauss_ds_1_update_0_stage_99;
      dark_weights_normed_gauss_ds_1_update_0_stage_101 <= dark_weights_normed_gauss_ds_1_update_0_stage_100;
      dark_weights_normed_gauss_ds_1_update_0_stage_102 <= dark_weights_normed_gauss_ds_1_update_0_stage_101;
      dark_weights_normed_gauss_ds_1_update_0_stage_103 <= dark_weights_normed_gauss_ds_1_update_0_stage_102;
      dark_weights_normed_gauss_ds_1_update_0_stage_104 <= dark_weights_normed_gauss_ds_1_update_0_stage_103;
      dark_weights_normed_gauss_ds_1_update_0_stage_105 <= dark_weights_normed_gauss_ds_1_update_0_stage_104;
      dark_weights_normed_gauss_ds_1_update_0_stage_106 <= dark_weights_normed_gauss_ds_1_update_0_stage_105;
      dark_weights_normed_gauss_ds_1_update_0_stage_107 <= dark_weights_normed_gauss_ds_1_update_0_stage_106;
      dark_weights_normed_gauss_ds_1_update_0_stage_108 <= dark_weights_normed_gauss_ds_1_update_0_stage_107;
      dark_weights_normed_gauss_ds_1_update_0_stage_109 <= dark_weights_normed_gauss_ds_1_update_0_stage_108;
      dark_weights_normed_gauss_ds_1_update_0_stage_110 <= dark_weights_normed_gauss_ds_1_update_0_stage_109;
      dark_weights_normed_gauss_ds_1_update_0_stage_111 <= dark_weights_normed_gauss_ds_1_update_0_stage_110;
      dark_weights_normed_gauss_ds_1_update_0_stage_112 <= dark_weights_normed_gauss_ds_1_update_0_stage_111;
      dark_weights_normed_gauss_ds_1_update_0_stage_113 <= dark_weights_normed_gauss_ds_1_update_0_stage_112;
      dark_weights_normed_gauss_ds_1_update_0_stage_114 <= dark_weights_normed_gauss_ds_1_update_0_stage_113;
      dark_weights_normed_gauss_ds_1_update_0_stage_115 <= dark_weights_normed_gauss_ds_1_update_0_stage_114;
      dark_weights_normed_gauss_ds_1_update_0_stage_116 <= dark_weights_normed_gauss_ds_1_update_0_stage_115;
      dark_weights_normed_gauss_ds_1_update_0_stage_117 <= dark_weights_normed_gauss_ds_1_update_0_stage_116;
      dark_weights_normed_gauss_ds_1_update_0_stage_118 <= dark_weights_normed_gauss_ds_1_update_0_stage_117;
      dark_weights_normed_gauss_ds_1_update_0_stage_119 <= dark_weights_normed_gauss_ds_1_update_0_stage_118;
      dark_weights_normed_gauss_ds_1_update_0_stage_120 <= dark_weights_normed_gauss_ds_1_update_0_stage_119;
      dark_weights_normed_gauss_ds_1_update_0_stage_121 <= dark_weights_normed_gauss_ds_1_update_0_stage_120;
      dark_weights_normed_gauss_ds_1_update_0_stage_122 <= dark_weights_normed_gauss_ds_1_update_0_stage_121;
      dark_weights_normed_gauss_ds_1_update_0_stage_123 <= dark_weights_normed_gauss_ds_1_update_0_stage_122;
      dark_weights_normed_gauss_ds_1_update_0_stage_124 <= dark_weights_normed_gauss_ds_1_update_0_stage_123;
      dark_weights_normed_gauss_ds_1_update_0_stage_125 <= dark_weights_normed_gauss_ds_1_update_0_stage_124;
      dark_weights_normed_gauss_ds_1_update_0_stage_126 <= dark_weights_normed_gauss_ds_1_update_0_stage_125;
      dark_weights_normed_gauss_ds_1_update_0_stage_127 <= dark_weights_normed_gauss_ds_1_update_0_stage_126;
      dark_weights_normed_gauss_ds_1_update_0_stage_128 <= dark_weights_normed_gauss_ds_1_update_0_stage_127;
      dark_weights_normed_gauss_ds_1_update_0_stage_129 <= dark_weights_normed_gauss_ds_1_update_0_stage_128;
      dark_weights_normed_gauss_ds_1_update_0_stage_130 <= dark_weights_normed_gauss_ds_1_update_0_stage_129;
      dark_weights_normed_gauss_ds_1_update_0_stage_131 <= dark_weights_normed_gauss_ds_1_update_0_stage_130;
      dark_weights_normed_gauss_ds_1_update_0_stage_132 <= dark_weights_normed_gauss_ds_1_update_0_stage_131;
      dark_weights_normed_gauss_ds_1_update_0_stage_133 <= dark_weights_normed_gauss_ds_1_update_0_stage_132;
      dark_weights_normed_gauss_ds_1_update_0_stage_134 <= dark_weights_normed_gauss_ds_1_update_0_stage_133;
      dark_weights_normed_gauss_ds_1_update_0_stage_135 <= dark_weights_normed_gauss_ds_1_update_0_stage_134;
      dark_weights_normed_gauss_ds_1_update_0_stage_136 <= dark_weights_normed_gauss_ds_1_update_0_stage_135;
      dark_weights_normed_gauss_ds_1_update_0_stage_137 <= dark_weights_normed_gauss_ds_1_update_0_stage_136;
      dark_weights_normed_gauss_ds_1_update_0_stage_138 <= dark_weights_normed_gauss_ds_1_update_0_stage_137;
      dark_weights_normed_gauss_ds_1_update_0_stage_139 <= dark_weights_normed_gauss_ds_1_update_0_stage_138;
      dark_weights_normed_gauss_ds_1_update_0_stage_140 <= dark_weights_normed_gauss_ds_1_update_0_stage_139;
      dark_weights_normed_gauss_ds_1_update_0_stage_141 <= dark_weights_normed_gauss_ds_1_update_0_stage_140;
      dark_weights_normed_gauss_ds_1_update_0_stage_142 <= dark_weights_normed_gauss_ds_1_update_0_stage_141;
      dark_weights_normed_gauss_ds_1_update_0_stage_143 <= dark_weights_normed_gauss_ds_1_update_0_stage_142;
      dark_weights_normed_gauss_ds_1_update_0_stage_144 <= dark_weights_normed_gauss_ds_1_update_0_stage_143;
      dark_weights_normed_gauss_ds_1_update_0_stage_145 <= dark_weights_normed_gauss_ds_1_update_0_stage_144;
      dark_weights_normed_gauss_ds_1_update_0_stage_146 <= dark_weights_normed_gauss_ds_1_update_0_stage_145;
      dark_weights_normed_gauss_ds_1_update_0_stage_147 <= dark_weights_normed_gauss_ds_1_update_0_stage_146;
      dark_weights_normed_gauss_ds_1_update_0_stage_148 <= dark_weights_normed_gauss_ds_1_update_0_stage_147;
      dark_weights_normed_gauss_ds_1_update_0_stage_149 <= dark_weights_normed_gauss_ds_1_update_0_stage_148;
      dark_weights_normed_gauss_ds_1_update_0_stage_150 <= dark_weights_normed_gauss_ds_1_update_0_stage_149;
      dark_weights_normed_gauss_ds_1_update_0_stage_151 <= dark_weights_normed_gauss_ds_1_update_0_stage_150;
      dark_weights_normed_gauss_ds_1_update_0_stage_152 <= dark_weights_normed_gauss_ds_1_update_0_stage_151;
      dark_weights_normed_gauss_ds_1_update_0_stage_153 <= dark_weights_normed_gauss_ds_1_update_0_stage_152;
      dark_weights_normed_gauss_ds_1_update_0_stage_154 <= dark_weights_normed_gauss_ds_1_update_0_stage_153;
      dark_weights_normed_gauss_ds_1_update_0_stage_155 <= dark_weights_normed_gauss_ds_1_update_0_stage_154;
      dark_weights_normed_gauss_ds_1_update_0_stage_156 <= dark_weights_normed_gauss_ds_1_update_0_stage_155;
      dark_weights_normed_gauss_ds_1_update_0_stage_157 <= dark_weights_normed_gauss_ds_1_update_0_stage_156;
      dark_weights_normed_gauss_ds_1_update_0_stage_158 <= dark_weights_normed_gauss_ds_1_update_0_stage_157;
      dark_weights_normed_gauss_ds_1_update_0_stage_159 <= dark_weights_normed_gauss_ds_1_update_0_stage_158;
      dark_weights_normed_gauss_ds_1_update_0_stage_160 <= dark_weights_normed_gauss_ds_1_update_0_stage_159;
      dark_weights_normed_gauss_ds_1_update_0_stage_161 <= dark_weights_normed_gauss_ds_1_update_0_stage_160;
      dark_weights_normed_gauss_ds_1_update_0_stage_162 <= dark_weights_normed_gauss_ds_1_update_0_stage_161;
      dark_weights_normed_gauss_ds_1_update_0_stage_163 <= dark_weights_normed_gauss_ds_1_update_0_stage_162;
      dark_weights_normed_gauss_ds_1_update_0_stage_164 <= dark_weights_normed_gauss_ds_1_update_0_stage_163;
      dark_weights_normed_gauss_ds_1_update_0_stage_165 <= dark_weights_normed_gauss_ds_1_update_0_stage_164;
      dark_weights_normed_gauss_ds_1_update_0_stage_166 <= dark_weights_normed_gauss_ds_1_update_0_stage_165;
      dark_weights_normed_gauss_ds_1_update_0_stage_167 <= dark_weights_normed_gauss_ds_1_update_0_stage_166;
      dark_weights_normed_gauss_ds_1_update_0_stage_168 <= dark_weights_normed_gauss_ds_1_update_0_stage_167;
      dark_weights_normed_gauss_ds_1_update_0_stage_169 <= dark_weights_normed_gauss_ds_1_update_0_stage_168;
      dark_weights_normed_gauss_ds_1_update_0_stage_170 <= dark_weights_normed_gauss_ds_1_update_0_stage_169;
      dark_weights_normed_gauss_ds_1_update_0_stage_171 <= dark_weights_normed_gauss_ds_1_update_0_stage_170;
      dark_weights_normed_gauss_ds_1_update_0_stage_172 <= dark_weights_normed_gauss_ds_1_update_0_stage_171;
      dark_weights_normed_gauss_ds_1_update_0_stage_173 <= dark_weights_normed_gauss_ds_1_update_0_stage_172;
      dark_weights_normed_gauss_ds_1_update_0_stage_174 <= dark_weights_normed_gauss_ds_1_update_0_stage_173;
      dark_weights_normed_gauss_ds_1_update_0_stage_175 <= dark_weights_normed_gauss_ds_1_update_0_stage_174;
      dark_weights_normed_gauss_ds_1_update_0_stage_176 <= dark_weights_normed_gauss_ds_1_update_0_stage_175;
      dark_weights_normed_gauss_ds_1_update_0_stage_177 <= dark_weights_normed_gauss_ds_1_update_0_stage_176;
      dark_weights_normed_gauss_ds_1_update_0_stage_178 <= dark_weights_normed_gauss_ds_1_update_0_stage_177;
      dark_weights_normed_gauss_ds_1_update_0_stage_179 <= dark_weights_normed_gauss_ds_1_update_0_stage_178;
      dark_weights_normed_gauss_ds_1_update_0_stage_180 <= dark_weights_normed_gauss_ds_1_update_0_stage_179;
      dark_weights_normed_gauss_ds_1_update_0_stage_181 <= dark_weights_normed_gauss_ds_1_update_0_stage_180;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_97 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_98 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_97;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_99 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_98;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_100 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_99;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_101 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_100;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_102 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_101;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_103 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_102;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_104 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_103;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_105 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_104;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_106 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_105;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_107 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_106;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_108 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_107;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_109 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_108;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_110 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_109;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_111 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_110;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_112 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_111;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_113 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_112;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_114 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_113;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_115 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_114;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_116 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_115;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_117 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_116;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_118 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_117;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_119 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_118;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_120 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_119;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_121 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_120;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_122 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_121;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_123 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_122;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_124 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_123;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_125 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_124;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_126 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_125;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_127 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_126;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_128 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_127;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_129 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_128;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_130 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_129;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_131 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_130;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_132 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_131;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_133 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_132;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_134 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_133;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_135 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_134;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_136 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_135;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_137 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_136;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_138 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_137;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_139 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_138;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_140 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_139;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_141 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_140;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_142 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_141;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_143 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_142;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_144 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_143;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_145 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_144;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_146 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_145;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_147 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_146;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_148 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_147;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_149 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_148;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_150 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_149;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_151 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_150;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_152 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_151;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_153 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_152;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_154 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_153;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_155 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_154;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_156 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_155;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_157 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_156;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_158 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_157;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_159 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_158;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_160 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_159;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_161 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_160;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_162 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_161;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_163 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_162;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_164 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_163;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_165 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_164;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_166 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_165;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_167 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_166;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_168 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_167;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_169 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_168;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_170 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_169;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_171 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_170;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_172 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_171;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_173 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_172;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_174 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_173;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_175 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_174;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_176 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_175;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_177 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_176;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_178 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_177;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_179 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_178;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_180 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_179;
      dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_181 <= dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65_stage_180;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_81 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_82 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_81;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_83 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_82;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_84 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_83;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_85 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_84;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_86 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_85;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_87 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_86;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_88 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_87;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_89 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_88;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_90 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_89;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_91 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_90;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_92 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_91;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_93 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_92;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_94 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_93;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_95 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_94;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_96 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_95;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_97 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_96;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_98 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_97;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_99 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_98;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_100 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_99;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_101 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_100;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_102 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_101;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_103 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_102;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_104 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_103;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_105 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_104;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_106 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_105;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_107 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_106;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_108 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_107;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_109 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_108;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_110 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_109;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_111 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_110;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_112 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_111;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_113 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_112;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_114 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_113;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_115 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_114;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_116 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_115;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_117 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_116;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_118 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_117;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_119 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_118;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_120 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_119;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_121 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_120;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_122 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_121;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_123 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_122;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_124 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_123;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_125 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_124;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_126 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_125;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_127 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_126;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_128 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_127;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_129 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_128;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_130 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_129;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_131 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_130;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_132 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_131;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_133 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_132;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_134 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_133;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_135 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_134;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_136 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_135;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_137 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_136;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_138 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_137;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_139 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_138;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_140 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_139;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_141 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_140;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_142 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_141;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_143 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_142;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_144 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_143;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_145 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_144;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_146 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_145;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_147 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_146;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_148 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_147;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_149 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_148;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_150 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_149;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_151 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_150;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_152 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_151;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_153 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_152;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_154 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_153;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_155 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_154;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_156 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_155;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_157 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_156;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_158 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_157;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_159 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_158;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_160 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_159;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_161 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_160;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_162 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_161;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_163 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_162;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_164 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_163;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_165 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_164;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_166 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_165;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_167 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_166;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_168 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_167;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_169 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_168;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_170 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_169;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_171 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_170;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_172 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_171;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_173 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_172;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_174 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_173;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_175 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_174;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_176 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_175;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_177 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_176;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_178 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_177;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_179 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_178;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_180 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_179;
      dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_181 <= dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54_stage_180;
      dark_gauss_blur_3_update_0_stage_98 <= dark_gauss_blur_3_update_0;
      dark_gauss_blur_3_update_0_stage_99 <= dark_gauss_blur_3_update_0_stage_98;
      dark_gauss_blur_3_update_0_stage_100 <= dark_gauss_blur_3_update_0_stage_99;
      dark_gauss_blur_3_update_0_stage_101 <= dark_gauss_blur_3_update_0_stage_100;
      dark_gauss_blur_3_update_0_stage_102 <= dark_gauss_blur_3_update_0_stage_101;
      dark_gauss_blur_3_update_0_stage_103 <= dark_gauss_blur_3_update_0_stage_102;
      dark_gauss_blur_3_update_0_stage_104 <= dark_gauss_blur_3_update_0_stage_103;
      dark_gauss_blur_3_update_0_stage_105 <= dark_gauss_blur_3_update_0_stage_104;
      dark_gauss_blur_3_update_0_stage_106 <= dark_gauss_blur_3_update_0_stage_105;
      dark_gauss_blur_3_update_0_stage_107 <= dark_gauss_blur_3_update_0_stage_106;
      dark_gauss_blur_3_update_0_stage_108 <= dark_gauss_blur_3_update_0_stage_107;
      dark_gauss_blur_3_update_0_stage_109 <= dark_gauss_blur_3_update_0_stage_108;
      dark_gauss_blur_3_update_0_stage_110 <= dark_gauss_blur_3_update_0_stage_109;
      dark_gauss_blur_3_update_0_stage_111 <= dark_gauss_blur_3_update_0_stage_110;
      dark_gauss_blur_3_update_0_stage_112 <= dark_gauss_blur_3_update_0_stage_111;
      dark_gauss_blur_3_update_0_stage_113 <= dark_gauss_blur_3_update_0_stage_112;
      dark_gauss_blur_3_update_0_stage_114 <= dark_gauss_blur_3_update_0_stage_113;
      dark_gauss_blur_3_update_0_stage_115 <= dark_gauss_blur_3_update_0_stage_114;
      dark_gauss_blur_3_update_0_stage_116 <= dark_gauss_blur_3_update_0_stage_115;
      dark_gauss_blur_3_update_0_stage_117 <= dark_gauss_blur_3_update_0_stage_116;
      dark_gauss_blur_3_update_0_stage_118 <= dark_gauss_blur_3_update_0_stage_117;
      dark_gauss_blur_3_update_0_stage_119 <= dark_gauss_blur_3_update_0_stage_118;
      dark_gauss_blur_3_update_0_stage_120 <= dark_gauss_blur_3_update_0_stage_119;
      dark_gauss_blur_3_update_0_stage_121 <= dark_gauss_blur_3_update_0_stage_120;
      dark_gauss_blur_3_update_0_stage_122 <= dark_gauss_blur_3_update_0_stage_121;
      dark_gauss_blur_3_update_0_stage_123 <= dark_gauss_blur_3_update_0_stage_122;
      dark_gauss_blur_3_update_0_stage_124 <= dark_gauss_blur_3_update_0_stage_123;
      dark_gauss_blur_3_update_0_stage_125 <= dark_gauss_blur_3_update_0_stage_124;
      dark_gauss_blur_3_update_0_stage_126 <= dark_gauss_blur_3_update_0_stage_125;
      dark_gauss_blur_3_update_0_stage_127 <= dark_gauss_blur_3_update_0_stage_126;
      dark_gauss_blur_3_update_0_stage_128 <= dark_gauss_blur_3_update_0_stage_127;
      dark_gauss_blur_3_update_0_stage_129 <= dark_gauss_blur_3_update_0_stage_128;
      dark_gauss_blur_3_update_0_stage_130 <= dark_gauss_blur_3_update_0_stage_129;
      dark_gauss_blur_3_update_0_stage_131 <= dark_gauss_blur_3_update_0_stage_130;
      dark_gauss_blur_3_update_0_stage_132 <= dark_gauss_blur_3_update_0_stage_131;
      dark_gauss_blur_3_update_0_stage_133 <= dark_gauss_blur_3_update_0_stage_132;
      dark_gauss_blur_3_update_0_stage_134 <= dark_gauss_blur_3_update_0_stage_133;
      dark_gauss_blur_3_update_0_stage_135 <= dark_gauss_blur_3_update_0_stage_134;
      dark_gauss_blur_3_update_0_stage_136 <= dark_gauss_blur_3_update_0_stage_135;
      dark_gauss_blur_3_update_0_stage_137 <= dark_gauss_blur_3_update_0_stage_136;
      dark_gauss_blur_3_update_0_stage_138 <= dark_gauss_blur_3_update_0_stage_137;
      dark_gauss_blur_3_update_0_stage_139 <= dark_gauss_blur_3_update_0_stage_138;
      dark_gauss_blur_3_update_0_stage_140 <= dark_gauss_blur_3_update_0_stage_139;
      dark_gauss_blur_3_update_0_stage_141 <= dark_gauss_blur_3_update_0_stage_140;
      dark_gauss_blur_3_update_0_stage_142 <= dark_gauss_blur_3_update_0_stage_141;
      dark_gauss_blur_3_update_0_stage_143 <= dark_gauss_blur_3_update_0_stage_142;
      dark_gauss_blur_3_update_0_stage_144 <= dark_gauss_blur_3_update_0_stage_143;
      dark_gauss_blur_3_update_0_stage_145 <= dark_gauss_blur_3_update_0_stage_144;
      dark_gauss_blur_3_update_0_stage_146 <= dark_gauss_blur_3_update_0_stage_145;
      dark_gauss_blur_3_update_0_stage_147 <= dark_gauss_blur_3_update_0_stage_146;
      dark_gauss_blur_3_update_0_stage_148 <= dark_gauss_blur_3_update_0_stage_147;
      dark_gauss_blur_3_update_0_stage_149 <= dark_gauss_blur_3_update_0_stage_148;
      dark_gauss_blur_3_update_0_stage_150 <= dark_gauss_blur_3_update_0_stage_149;
      dark_gauss_blur_3_update_0_stage_151 <= dark_gauss_blur_3_update_0_stage_150;
      dark_gauss_blur_3_update_0_stage_152 <= dark_gauss_blur_3_update_0_stage_151;
      dark_gauss_blur_3_update_0_stage_153 <= dark_gauss_blur_3_update_0_stage_152;
      dark_gauss_blur_3_update_0_stage_154 <= dark_gauss_blur_3_update_0_stage_153;
      dark_gauss_blur_3_update_0_stage_155 <= dark_gauss_blur_3_update_0_stage_154;
      dark_gauss_blur_3_update_0_stage_156 <= dark_gauss_blur_3_update_0_stage_155;
      dark_gauss_blur_3_update_0_stage_157 <= dark_gauss_blur_3_update_0_stage_156;
      dark_gauss_blur_3_update_0_stage_158 <= dark_gauss_blur_3_update_0_stage_157;
      dark_gauss_blur_3_update_0_stage_159 <= dark_gauss_blur_3_update_0_stage_158;
      dark_gauss_blur_3_update_0_stage_160 <= dark_gauss_blur_3_update_0_stage_159;
      dark_gauss_blur_3_update_0_stage_161 <= dark_gauss_blur_3_update_0_stage_160;
      dark_gauss_blur_3_update_0_stage_162 <= dark_gauss_blur_3_update_0_stage_161;
      dark_gauss_blur_3_update_0_stage_163 <= dark_gauss_blur_3_update_0_stage_162;
      dark_gauss_blur_3_update_0_stage_164 <= dark_gauss_blur_3_update_0_stage_163;
      dark_gauss_blur_3_update_0_stage_165 <= dark_gauss_blur_3_update_0_stage_164;
      dark_gauss_blur_3_update_0_stage_166 <= dark_gauss_blur_3_update_0_stage_165;
      dark_gauss_blur_3_update_0_stage_167 <= dark_gauss_blur_3_update_0_stage_166;
      dark_gauss_blur_3_update_0_stage_168 <= dark_gauss_blur_3_update_0_stage_167;
      dark_gauss_blur_3_update_0_stage_169 <= dark_gauss_blur_3_update_0_stage_168;
      dark_gauss_blur_3_update_0_stage_170 <= dark_gauss_blur_3_update_0_stage_169;
      dark_gauss_blur_3_update_0_stage_171 <= dark_gauss_blur_3_update_0_stage_170;
      dark_gauss_blur_3_update_0_stage_172 <= dark_gauss_blur_3_update_0_stage_171;
      dark_gauss_blur_3_update_0_stage_173 <= dark_gauss_blur_3_update_0_stage_172;
      dark_gauss_blur_3_update_0_stage_174 <= dark_gauss_blur_3_update_0_stage_173;
      dark_gauss_blur_3_update_0_stage_175 <= dark_gauss_blur_3_update_0_stage_174;
      dark_gauss_blur_3_update_0_stage_176 <= dark_gauss_blur_3_update_0_stage_175;
      dark_gauss_blur_3_update_0_stage_177 <= dark_gauss_blur_3_update_0_stage_176;
      dark_gauss_blur_3_update_0_stage_178 <= dark_gauss_blur_3_update_0_stage_177;
      dark_gauss_blur_3_update_0_stage_179 <= dark_gauss_blur_3_update_0_stage_178;
      dark_gauss_blur_3_update_0_stage_180 <= dark_gauss_blur_3_update_0_stage_179;
      dark_gauss_blur_3_update_0_stage_181 <= dark_gauss_blur_3_update_0_stage_180;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_99 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_100 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_99;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_101 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_100;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_102 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_101;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_103 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_102;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_104 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_103;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_105 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_104;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_106 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_105;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_107 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_106;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_108 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_107;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_109 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_108;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_110 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_109;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_111 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_110;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_112 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_111;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_113 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_112;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_114 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_113;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_115 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_114;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_116 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_115;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_117 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_116;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_118 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_117;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_119 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_118;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_120 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_119;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_121 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_120;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_122 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_121;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_123 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_122;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_124 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_123;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_125 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_124;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_126 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_125;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_127 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_126;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_128 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_127;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_129 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_128;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_130 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_129;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_131 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_130;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_132 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_131;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_133 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_132;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_134 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_133;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_135 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_134;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_136 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_135;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_137 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_136;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_138 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_137;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_139 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_138;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_140 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_139;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_141 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_140;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_142 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_141;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_143 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_142;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_144 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_143;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_145 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_144;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_146 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_145;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_147 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_146;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_148 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_147;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_149 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_148;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_150 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_149;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_151 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_150;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_152 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_151;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_153 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_152;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_154 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_153;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_155 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_154;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_156 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_155;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_157 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_156;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_158 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_157;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_159 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_158;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_160 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_159;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_161 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_160;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_162 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_161;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_163 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_162;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_164 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_163;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_165 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_164;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_166 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_165;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_167 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_166;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_168 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_167;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_169 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_168;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_170 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_169;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_171 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_170;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_172 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_171;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_173 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_172;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_174 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_173;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_175 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_174;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_176 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_175;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_177 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_176;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_178 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_177;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_179 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_178;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_180 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_179;
      dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_181 <= dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66_stage_180;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_104 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_105 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_104;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_106 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_105;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_107 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_106;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_108 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_107;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_109 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_108;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_110 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_109;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_111 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_110;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_112 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_111;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_113 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_112;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_114 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_113;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_115 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_114;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_116 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_115;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_117 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_116;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_118 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_117;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_119 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_118;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_120 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_119;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_121 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_120;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_122 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_121;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_123 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_122;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_124 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_123;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_125 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_124;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_126 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_125;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_127 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_126;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_128 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_127;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_129 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_128;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_130 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_129;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_131 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_130;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_132 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_131;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_133 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_132;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_134 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_133;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_135 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_134;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_136 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_135;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_137 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_136;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_138 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_137;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_139 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_138;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_140 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_139;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_141 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_140;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_142 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_141;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_143 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_142;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_144 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_143;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_145 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_144;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_146 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_145;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_147 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_146;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_148 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_147;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_149 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_148;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_150 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_149;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_151 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_150;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_152 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_151;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_153 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_152;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_154 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_153;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_155 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_154;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_156 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_155;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_157 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_156;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_158 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_157;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_159 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_158;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_160 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_159;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_161 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_160;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_162 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_161;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_163 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_162;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_164 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_163;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_165 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_164;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_166 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_165;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_167 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_166;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_168 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_167;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_169 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_168;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_170 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_169;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_171 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_170;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_172 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_171;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_173 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_172;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_174 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_173;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_175 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_174;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_176 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_175;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_177 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_176;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_178 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_177;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_179 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_178;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_180 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_179;
      bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_181 <= bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70_stage_180;
      bright_weights_normed_gauss_ds_1_update_0_stage_105 <= bright_weights_normed_gauss_ds_1_update_0;
      bright_weights_normed_gauss_ds_1_update_0_stage_106 <= bright_weights_normed_gauss_ds_1_update_0_stage_105;
      bright_weights_normed_gauss_ds_1_update_0_stage_107 <= bright_weights_normed_gauss_ds_1_update_0_stage_106;
      bright_weights_normed_gauss_ds_1_update_0_stage_108 <= bright_weights_normed_gauss_ds_1_update_0_stage_107;
      bright_weights_normed_gauss_ds_1_update_0_stage_109 <= bright_weights_normed_gauss_ds_1_update_0_stage_108;
      bright_weights_normed_gauss_ds_1_update_0_stage_110 <= bright_weights_normed_gauss_ds_1_update_0_stage_109;
      bright_weights_normed_gauss_ds_1_update_0_stage_111 <= bright_weights_normed_gauss_ds_1_update_0_stage_110;
      bright_weights_normed_gauss_ds_1_update_0_stage_112 <= bright_weights_normed_gauss_ds_1_update_0_stage_111;
      bright_weights_normed_gauss_ds_1_update_0_stage_113 <= bright_weights_normed_gauss_ds_1_update_0_stage_112;
      bright_weights_normed_gauss_ds_1_update_0_stage_114 <= bright_weights_normed_gauss_ds_1_update_0_stage_113;
      bright_weights_normed_gauss_ds_1_update_0_stage_115 <= bright_weights_normed_gauss_ds_1_update_0_stage_114;
      bright_weights_normed_gauss_ds_1_update_0_stage_116 <= bright_weights_normed_gauss_ds_1_update_0_stage_115;
      bright_weights_normed_gauss_ds_1_update_0_stage_117 <= bright_weights_normed_gauss_ds_1_update_0_stage_116;
      bright_weights_normed_gauss_ds_1_update_0_stage_118 <= bright_weights_normed_gauss_ds_1_update_0_stage_117;
      bright_weights_normed_gauss_ds_1_update_0_stage_119 <= bright_weights_normed_gauss_ds_1_update_0_stage_118;
      bright_weights_normed_gauss_ds_1_update_0_stage_120 <= bright_weights_normed_gauss_ds_1_update_0_stage_119;
      bright_weights_normed_gauss_ds_1_update_0_stage_121 <= bright_weights_normed_gauss_ds_1_update_0_stage_120;
      bright_weights_normed_gauss_ds_1_update_0_stage_122 <= bright_weights_normed_gauss_ds_1_update_0_stage_121;
      bright_weights_normed_gauss_ds_1_update_0_stage_123 <= bright_weights_normed_gauss_ds_1_update_0_stage_122;
      bright_weights_normed_gauss_ds_1_update_0_stage_124 <= bright_weights_normed_gauss_ds_1_update_0_stage_123;
      bright_weights_normed_gauss_ds_1_update_0_stage_125 <= bright_weights_normed_gauss_ds_1_update_0_stage_124;
      bright_weights_normed_gauss_ds_1_update_0_stage_126 <= bright_weights_normed_gauss_ds_1_update_0_stage_125;
      bright_weights_normed_gauss_ds_1_update_0_stage_127 <= bright_weights_normed_gauss_ds_1_update_0_stage_126;
      bright_weights_normed_gauss_ds_1_update_0_stage_128 <= bright_weights_normed_gauss_ds_1_update_0_stage_127;
      bright_weights_normed_gauss_ds_1_update_0_stage_129 <= bright_weights_normed_gauss_ds_1_update_0_stage_128;
      bright_weights_normed_gauss_ds_1_update_0_stage_130 <= bright_weights_normed_gauss_ds_1_update_0_stage_129;
      bright_weights_normed_gauss_ds_1_update_0_stage_131 <= bright_weights_normed_gauss_ds_1_update_0_stage_130;
      bright_weights_normed_gauss_ds_1_update_0_stage_132 <= bright_weights_normed_gauss_ds_1_update_0_stage_131;
      bright_weights_normed_gauss_ds_1_update_0_stage_133 <= bright_weights_normed_gauss_ds_1_update_0_stage_132;
      bright_weights_normed_gauss_ds_1_update_0_stage_134 <= bright_weights_normed_gauss_ds_1_update_0_stage_133;
      bright_weights_normed_gauss_ds_1_update_0_stage_135 <= bright_weights_normed_gauss_ds_1_update_0_stage_134;
      bright_weights_normed_gauss_ds_1_update_0_stage_136 <= bright_weights_normed_gauss_ds_1_update_0_stage_135;
      bright_weights_normed_gauss_ds_1_update_0_stage_137 <= bright_weights_normed_gauss_ds_1_update_0_stage_136;
      bright_weights_normed_gauss_ds_1_update_0_stage_138 <= bright_weights_normed_gauss_ds_1_update_0_stage_137;
      bright_weights_normed_gauss_ds_1_update_0_stage_139 <= bright_weights_normed_gauss_ds_1_update_0_stage_138;
      bright_weights_normed_gauss_ds_1_update_0_stage_140 <= bright_weights_normed_gauss_ds_1_update_0_stage_139;
      bright_weights_normed_gauss_ds_1_update_0_stage_141 <= bright_weights_normed_gauss_ds_1_update_0_stage_140;
      bright_weights_normed_gauss_ds_1_update_0_stage_142 <= bright_weights_normed_gauss_ds_1_update_0_stage_141;
      bright_weights_normed_gauss_ds_1_update_0_stage_143 <= bright_weights_normed_gauss_ds_1_update_0_stage_142;
      bright_weights_normed_gauss_ds_1_update_0_stage_144 <= bright_weights_normed_gauss_ds_1_update_0_stage_143;
      bright_weights_normed_gauss_ds_1_update_0_stage_145 <= bright_weights_normed_gauss_ds_1_update_0_stage_144;
      bright_weights_normed_gauss_ds_1_update_0_stage_146 <= bright_weights_normed_gauss_ds_1_update_0_stage_145;
      bright_weights_normed_gauss_ds_1_update_0_stage_147 <= bright_weights_normed_gauss_ds_1_update_0_stage_146;
      bright_weights_normed_gauss_ds_1_update_0_stage_148 <= bright_weights_normed_gauss_ds_1_update_0_stage_147;
      bright_weights_normed_gauss_ds_1_update_0_stage_149 <= bright_weights_normed_gauss_ds_1_update_0_stage_148;
      bright_weights_normed_gauss_ds_1_update_0_stage_150 <= bright_weights_normed_gauss_ds_1_update_0_stage_149;
      bright_weights_normed_gauss_ds_1_update_0_stage_151 <= bright_weights_normed_gauss_ds_1_update_0_stage_150;
      bright_weights_normed_gauss_ds_1_update_0_stage_152 <= bright_weights_normed_gauss_ds_1_update_0_stage_151;
      bright_weights_normed_gauss_ds_1_update_0_stage_153 <= bright_weights_normed_gauss_ds_1_update_0_stage_152;
      bright_weights_normed_gauss_ds_1_update_0_stage_154 <= bright_weights_normed_gauss_ds_1_update_0_stage_153;
      bright_weights_normed_gauss_ds_1_update_0_stage_155 <= bright_weights_normed_gauss_ds_1_update_0_stage_154;
      bright_weights_normed_gauss_ds_1_update_0_stage_156 <= bright_weights_normed_gauss_ds_1_update_0_stage_155;
      bright_weights_normed_gauss_ds_1_update_0_stage_157 <= bright_weights_normed_gauss_ds_1_update_0_stage_156;
      bright_weights_normed_gauss_ds_1_update_0_stage_158 <= bright_weights_normed_gauss_ds_1_update_0_stage_157;
      bright_weights_normed_gauss_ds_1_update_0_stage_159 <= bright_weights_normed_gauss_ds_1_update_0_stage_158;
      bright_weights_normed_gauss_ds_1_update_0_stage_160 <= bright_weights_normed_gauss_ds_1_update_0_stage_159;
      bright_weights_normed_gauss_ds_1_update_0_stage_161 <= bright_weights_normed_gauss_ds_1_update_0_stage_160;
      bright_weights_normed_gauss_ds_1_update_0_stage_162 <= bright_weights_normed_gauss_ds_1_update_0_stage_161;
      bright_weights_normed_gauss_ds_1_update_0_stage_163 <= bright_weights_normed_gauss_ds_1_update_0_stage_162;
      bright_weights_normed_gauss_ds_1_update_0_stage_164 <= bright_weights_normed_gauss_ds_1_update_0_stage_163;
      bright_weights_normed_gauss_ds_1_update_0_stage_165 <= bright_weights_normed_gauss_ds_1_update_0_stage_164;
      bright_weights_normed_gauss_ds_1_update_0_stage_166 <= bright_weights_normed_gauss_ds_1_update_0_stage_165;
      bright_weights_normed_gauss_ds_1_update_0_stage_167 <= bright_weights_normed_gauss_ds_1_update_0_stage_166;
      bright_weights_normed_gauss_ds_1_update_0_stage_168 <= bright_weights_normed_gauss_ds_1_update_0_stage_167;
      bright_weights_normed_gauss_ds_1_update_0_stage_169 <= bright_weights_normed_gauss_ds_1_update_0_stage_168;
      bright_weights_normed_gauss_ds_1_update_0_stage_170 <= bright_weights_normed_gauss_ds_1_update_0_stage_169;
      bright_weights_normed_gauss_ds_1_update_0_stage_171 <= bright_weights_normed_gauss_ds_1_update_0_stage_170;
      bright_weights_normed_gauss_ds_1_update_0_stage_172 <= bright_weights_normed_gauss_ds_1_update_0_stage_171;
      bright_weights_normed_gauss_ds_1_update_0_stage_173 <= bright_weights_normed_gauss_ds_1_update_0_stage_172;
      bright_weights_normed_gauss_ds_1_update_0_stage_174 <= bright_weights_normed_gauss_ds_1_update_0_stage_173;
      bright_weights_normed_gauss_ds_1_update_0_stage_175 <= bright_weights_normed_gauss_ds_1_update_0_stage_174;
      bright_weights_normed_gauss_ds_1_update_0_stage_176 <= bright_weights_normed_gauss_ds_1_update_0_stage_175;
      bright_weights_normed_gauss_ds_1_update_0_stage_177 <= bright_weights_normed_gauss_ds_1_update_0_stage_176;
      bright_weights_normed_gauss_ds_1_update_0_stage_178 <= bright_weights_normed_gauss_ds_1_update_0_stage_177;
      bright_weights_normed_gauss_ds_1_update_0_stage_179 <= bright_weights_normed_gauss_ds_1_update_0_stage_178;
      bright_weights_normed_gauss_ds_1_update_0_stage_180 <= bright_weights_normed_gauss_ds_1_update_0_stage_179;
      bright_weights_normed_gauss_ds_1_update_0_stage_181 <= bright_weights_normed_gauss_ds_1_update_0_stage_180;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_106 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_107 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_106;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_108 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_107;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_109 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_108;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_110 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_109;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_111 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_110;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_112 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_111;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_113 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_112;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_114 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_113;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_115 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_114;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_116 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_115;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_117 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_116;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_118 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_117;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_119 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_118;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_120 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_119;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_121 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_120;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_122 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_121;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_123 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_122;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_124 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_123;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_125 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_124;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_126 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_125;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_127 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_126;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_128 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_127;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_129 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_128;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_130 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_129;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_131 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_130;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_132 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_131;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_133 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_132;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_134 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_133;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_135 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_134;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_136 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_135;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_137 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_136;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_138 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_137;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_139 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_138;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_140 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_139;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_141 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_140;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_142 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_141;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_143 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_142;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_144 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_143;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_145 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_144;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_146 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_145;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_147 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_146;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_148 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_147;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_149 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_148;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_150 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_149;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_151 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_150;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_152 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_151;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_153 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_152;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_154 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_153;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_155 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_154;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_156 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_155;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_157 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_156;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_158 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_157;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_159 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_158;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_160 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_159;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_161 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_160;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_162 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_161;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_163 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_162;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_164 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_163;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_165 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_164;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_166 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_165;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_167 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_166;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_168 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_167;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_169 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_168;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_170 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_169;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_171 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_170;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_172 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_171;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_173 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_172;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_174 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_173;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_175 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_174;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_176 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_175;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_177 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_176;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_178 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_177;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_179 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_178;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_180 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_179;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_181 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71_stage_180;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_126 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_127 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_126;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_128 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_127;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_129 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_128;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_130 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_129;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_131 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_130;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_132 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_131;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_133 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_132;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_134 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_133;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_135 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_134;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_136 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_135;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_137 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_136;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_138 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_137;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_139 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_138;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_140 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_139;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_141 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_140;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_142 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_141;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_143 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_142;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_144 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_143;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_145 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_144;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_146 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_145;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_147 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_146;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_148 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_147;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_149 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_148;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_150 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_149;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_151 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_150;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_152 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_151;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_153 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_152;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_154 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_153;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_155 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_154;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_156 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_155;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_157 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_156;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_158 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_157;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_159 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_158;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_160 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_159;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_161 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_160;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_162 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_161;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_163 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_162;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_164 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_163;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_165 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_164;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_166 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_165;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_167 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_166;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_168 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_167;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_169 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_168;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_170 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_169;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_171 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_170;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_172 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_171;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_173 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_172;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_174 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_173;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_175 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_174;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_176 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_175;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_177 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_176;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_178 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_177;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_179 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_178;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_180 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_179;
      bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_181 <= bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87_stage_180;
      fused_level_1_update_0_stage_128 <= fused_level_1_update_0;
      fused_level_1_update_0_stage_129 <= fused_level_1_update_0_stage_128;
      fused_level_1_update_0_stage_130 <= fused_level_1_update_0_stage_129;
      fused_level_1_update_0_stage_131 <= fused_level_1_update_0_stage_130;
      fused_level_1_update_0_stage_132 <= fused_level_1_update_0_stage_131;
      fused_level_1_update_0_stage_133 <= fused_level_1_update_0_stage_132;
      fused_level_1_update_0_stage_134 <= fused_level_1_update_0_stage_133;
      fused_level_1_update_0_stage_135 <= fused_level_1_update_0_stage_134;
      fused_level_1_update_0_stage_136 <= fused_level_1_update_0_stage_135;
      fused_level_1_update_0_stage_137 <= fused_level_1_update_0_stage_136;
      fused_level_1_update_0_stage_138 <= fused_level_1_update_0_stage_137;
      fused_level_1_update_0_stage_139 <= fused_level_1_update_0_stage_138;
      fused_level_1_update_0_stage_140 <= fused_level_1_update_0_stage_139;
      fused_level_1_update_0_stage_141 <= fused_level_1_update_0_stage_140;
      fused_level_1_update_0_stage_142 <= fused_level_1_update_0_stage_141;
      fused_level_1_update_0_stage_143 <= fused_level_1_update_0_stage_142;
      fused_level_1_update_0_stage_144 <= fused_level_1_update_0_stage_143;
      fused_level_1_update_0_stage_145 <= fused_level_1_update_0_stage_144;
      fused_level_1_update_0_stage_146 <= fused_level_1_update_0_stage_145;
      fused_level_1_update_0_stage_147 <= fused_level_1_update_0_stage_146;
      fused_level_1_update_0_stage_148 <= fused_level_1_update_0_stage_147;
      fused_level_1_update_0_stage_149 <= fused_level_1_update_0_stage_148;
      fused_level_1_update_0_stage_150 <= fused_level_1_update_0_stage_149;
      fused_level_1_update_0_stage_151 <= fused_level_1_update_0_stage_150;
      fused_level_1_update_0_stage_152 <= fused_level_1_update_0_stage_151;
      fused_level_1_update_0_stage_153 <= fused_level_1_update_0_stage_152;
      fused_level_1_update_0_stage_154 <= fused_level_1_update_0_stage_153;
      fused_level_1_update_0_stage_155 <= fused_level_1_update_0_stage_154;
      fused_level_1_update_0_stage_156 <= fused_level_1_update_0_stage_155;
      fused_level_1_update_0_stage_157 <= fused_level_1_update_0_stage_156;
      fused_level_1_update_0_stage_158 <= fused_level_1_update_0_stage_157;
      fused_level_1_update_0_stage_159 <= fused_level_1_update_0_stage_158;
      fused_level_1_update_0_stage_160 <= fused_level_1_update_0_stage_159;
      fused_level_1_update_0_stage_161 <= fused_level_1_update_0_stage_160;
      fused_level_1_update_0_stage_162 <= fused_level_1_update_0_stage_161;
      fused_level_1_update_0_stage_163 <= fused_level_1_update_0_stage_162;
      fused_level_1_update_0_stage_164 <= fused_level_1_update_0_stage_163;
      fused_level_1_update_0_stage_165 <= fused_level_1_update_0_stage_164;
      fused_level_1_update_0_stage_166 <= fused_level_1_update_0_stage_165;
      fused_level_1_update_0_stage_167 <= fused_level_1_update_0_stage_166;
      fused_level_1_update_0_stage_168 <= fused_level_1_update_0_stage_167;
      fused_level_1_update_0_stage_169 <= fused_level_1_update_0_stage_168;
      fused_level_1_update_0_stage_170 <= fused_level_1_update_0_stage_169;
      fused_level_1_update_0_stage_171 <= fused_level_1_update_0_stage_170;
      fused_level_1_update_0_stage_172 <= fused_level_1_update_0_stage_171;
      fused_level_1_update_0_stage_173 <= fused_level_1_update_0_stage_172;
      fused_level_1_update_0_stage_174 <= fused_level_1_update_0_stage_173;
      fused_level_1_update_0_stage_175 <= fused_level_1_update_0_stage_174;
      fused_level_1_update_0_stage_176 <= fused_level_1_update_0_stage_175;
      fused_level_1_update_0_stage_177 <= fused_level_1_update_0_stage_176;
      fused_level_1_update_0_stage_178 <= fused_level_1_update_0_stage_177;
      fused_level_1_update_0_stage_179 <= fused_level_1_update_0_stage_178;
      fused_level_1_update_0_stage_180 <= fused_level_1_update_0_stage_179;
      fused_level_1_update_0_stage_181 <= fused_level_1_update_0_stage_180;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_127 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_128 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_127;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_129 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_128;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_130 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_129;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_131 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_130;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_132 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_131;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_133 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_132;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_134 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_133;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_135 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_134;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_136 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_135;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_137 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_136;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_138 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_137;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_139 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_138;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_140 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_139;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_141 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_140;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_142 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_141;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_143 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_142;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_144 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_143;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_145 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_144;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_146 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_145;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_147 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_146;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_148 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_147;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_149 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_148;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_150 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_149;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_151 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_150;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_152 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_151;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_153 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_152;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_154 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_153;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_155 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_154;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_156 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_155;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_157 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_156;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_158 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_157;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_159 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_158;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_160 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_159;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_161 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_160;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_162 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_161;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_163 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_162;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_164 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_163;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_165 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_164;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_166 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_165;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_167 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_166;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_168 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_167;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_169 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_168;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_170 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_169;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_171 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_170;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_172 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_171;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_173 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_172;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_174 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_173;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_175 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_174;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_176 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_175;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_177 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_176;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_178 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_177;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_179 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_178;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_180 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_179;
      dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_181 <= dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88_stage_180;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_129 <= fused_level_1_fused_level_1_update_0_write_write_89;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_130 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_129;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_131 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_130;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_132 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_131;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_133 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_132;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_134 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_133;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_135 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_134;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_136 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_135;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_137 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_136;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_138 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_137;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_139 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_138;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_140 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_139;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_141 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_140;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_142 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_141;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_143 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_142;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_144 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_143;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_145 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_144;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_146 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_145;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_147 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_146;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_148 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_147;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_149 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_148;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_150 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_149;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_151 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_150;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_152 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_151;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_153 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_152;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_154 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_153;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_155 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_154;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_156 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_155;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_157 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_156;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_158 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_157;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_159 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_158;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_160 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_159;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_161 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_160;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_162 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_161;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_163 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_162;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_164 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_163;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_165 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_164;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_166 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_165;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_167 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_166;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_168 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_167;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_169 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_168;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_170 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_169;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_171 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_170;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_172 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_171;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_173 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_172;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_174 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_173;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_175 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_174;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_176 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_175;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_177 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_176;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_178 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_177;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_179 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_178;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_180 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_179;
      fused_level_1_fused_level_1_update_0_write_write_89_stage_181 <= fused_level_1_fused_level_1_update_0_write_write_89_stage_180;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_136 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_137 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_136;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_138 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_137;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_139 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_138;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_140 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_139;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_141 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_140;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_142 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_141;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_143 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_142;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_144 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_143;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_145 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_144;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_146 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_145;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_147 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_146;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_148 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_147;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_149 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_148;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_150 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_149;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_151 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_150;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_152 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_151;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_153 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_152;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_154 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_153;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_155 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_154;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_156 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_155;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_157 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_156;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_158 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_157;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_159 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_158;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_160 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_159;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_161 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_160;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_162 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_161;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_163 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_162;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_164 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_163;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_165 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_164;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_166 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_165;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_167 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_166;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_168 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_167;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_169 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_168;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_170 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_169;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_171 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_170;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_172 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_171;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_173 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_172;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_174 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_173;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_175 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_174;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_176 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_175;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_177 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_176;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_178 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_177;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_179 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_178;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_180 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_179;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_181 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94_stage_180;
      dark_weights_normed_gauss_ds_3_update_0_stage_137 <= dark_weights_normed_gauss_ds_3_update_0;
      dark_weights_normed_gauss_ds_3_update_0_stage_138 <= dark_weights_normed_gauss_ds_3_update_0_stage_137;
      dark_weights_normed_gauss_ds_3_update_0_stage_139 <= dark_weights_normed_gauss_ds_3_update_0_stage_138;
      dark_weights_normed_gauss_ds_3_update_0_stage_140 <= dark_weights_normed_gauss_ds_3_update_0_stage_139;
      dark_weights_normed_gauss_ds_3_update_0_stage_141 <= dark_weights_normed_gauss_ds_3_update_0_stage_140;
      dark_weights_normed_gauss_ds_3_update_0_stage_142 <= dark_weights_normed_gauss_ds_3_update_0_stage_141;
      dark_weights_normed_gauss_ds_3_update_0_stage_143 <= dark_weights_normed_gauss_ds_3_update_0_stage_142;
      dark_weights_normed_gauss_ds_3_update_0_stage_144 <= dark_weights_normed_gauss_ds_3_update_0_stage_143;
      dark_weights_normed_gauss_ds_3_update_0_stage_145 <= dark_weights_normed_gauss_ds_3_update_0_stage_144;
      dark_weights_normed_gauss_ds_3_update_0_stage_146 <= dark_weights_normed_gauss_ds_3_update_0_stage_145;
      dark_weights_normed_gauss_ds_3_update_0_stage_147 <= dark_weights_normed_gauss_ds_3_update_0_stage_146;
      dark_weights_normed_gauss_ds_3_update_0_stage_148 <= dark_weights_normed_gauss_ds_3_update_0_stage_147;
      dark_weights_normed_gauss_ds_3_update_0_stage_149 <= dark_weights_normed_gauss_ds_3_update_0_stage_148;
      dark_weights_normed_gauss_ds_3_update_0_stage_150 <= dark_weights_normed_gauss_ds_3_update_0_stage_149;
      dark_weights_normed_gauss_ds_3_update_0_stage_151 <= dark_weights_normed_gauss_ds_3_update_0_stage_150;
      dark_weights_normed_gauss_ds_3_update_0_stage_152 <= dark_weights_normed_gauss_ds_3_update_0_stage_151;
      dark_weights_normed_gauss_ds_3_update_0_stage_153 <= dark_weights_normed_gauss_ds_3_update_0_stage_152;
      dark_weights_normed_gauss_ds_3_update_0_stage_154 <= dark_weights_normed_gauss_ds_3_update_0_stage_153;
      dark_weights_normed_gauss_ds_3_update_0_stage_155 <= dark_weights_normed_gauss_ds_3_update_0_stage_154;
      dark_weights_normed_gauss_ds_3_update_0_stage_156 <= dark_weights_normed_gauss_ds_3_update_0_stage_155;
      dark_weights_normed_gauss_ds_3_update_0_stage_157 <= dark_weights_normed_gauss_ds_3_update_0_stage_156;
      dark_weights_normed_gauss_ds_3_update_0_stage_158 <= dark_weights_normed_gauss_ds_3_update_0_stage_157;
      dark_weights_normed_gauss_ds_3_update_0_stage_159 <= dark_weights_normed_gauss_ds_3_update_0_stage_158;
      dark_weights_normed_gauss_ds_3_update_0_stage_160 <= dark_weights_normed_gauss_ds_3_update_0_stage_159;
      dark_weights_normed_gauss_ds_3_update_0_stage_161 <= dark_weights_normed_gauss_ds_3_update_0_stage_160;
      dark_weights_normed_gauss_ds_3_update_0_stage_162 <= dark_weights_normed_gauss_ds_3_update_0_stage_161;
      dark_weights_normed_gauss_ds_3_update_0_stage_163 <= dark_weights_normed_gauss_ds_3_update_0_stage_162;
      dark_weights_normed_gauss_ds_3_update_0_stage_164 <= dark_weights_normed_gauss_ds_3_update_0_stage_163;
      dark_weights_normed_gauss_ds_3_update_0_stage_165 <= dark_weights_normed_gauss_ds_3_update_0_stage_164;
      dark_weights_normed_gauss_ds_3_update_0_stage_166 <= dark_weights_normed_gauss_ds_3_update_0_stage_165;
      dark_weights_normed_gauss_ds_3_update_0_stage_167 <= dark_weights_normed_gauss_ds_3_update_0_stage_166;
      dark_weights_normed_gauss_ds_3_update_0_stage_168 <= dark_weights_normed_gauss_ds_3_update_0_stage_167;
      dark_weights_normed_gauss_ds_3_update_0_stage_169 <= dark_weights_normed_gauss_ds_3_update_0_stage_168;
      dark_weights_normed_gauss_ds_3_update_0_stage_170 <= dark_weights_normed_gauss_ds_3_update_0_stage_169;
      dark_weights_normed_gauss_ds_3_update_0_stage_171 <= dark_weights_normed_gauss_ds_3_update_0_stage_170;
      dark_weights_normed_gauss_ds_3_update_0_stage_172 <= dark_weights_normed_gauss_ds_3_update_0_stage_171;
      dark_weights_normed_gauss_ds_3_update_0_stage_173 <= dark_weights_normed_gauss_ds_3_update_0_stage_172;
      dark_weights_normed_gauss_ds_3_update_0_stage_174 <= dark_weights_normed_gauss_ds_3_update_0_stage_173;
      dark_weights_normed_gauss_ds_3_update_0_stage_175 <= dark_weights_normed_gauss_ds_3_update_0_stage_174;
      dark_weights_normed_gauss_ds_3_update_0_stage_176 <= dark_weights_normed_gauss_ds_3_update_0_stage_175;
      dark_weights_normed_gauss_ds_3_update_0_stage_177 <= dark_weights_normed_gauss_ds_3_update_0_stage_176;
      dark_weights_normed_gauss_ds_3_update_0_stage_178 <= dark_weights_normed_gauss_ds_3_update_0_stage_177;
      dark_weights_normed_gauss_ds_3_update_0_stage_179 <= dark_weights_normed_gauss_ds_3_update_0_stage_178;
      dark_weights_normed_gauss_ds_3_update_0_stage_180 <= dark_weights_normed_gauss_ds_3_update_0_stage_179;
      dark_weights_normed_gauss_ds_3_update_0_stage_181 <= dark_weights_normed_gauss_ds_3_update_0_stage_180;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_142 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_143 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_142;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_144 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_143;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_145 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_144;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_146 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_145;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_147 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_146;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_148 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_147;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_149 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_148;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_150 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_149;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_151 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_150;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_152 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_151;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_153 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_152;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_154 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_153;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_155 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_154;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_156 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_155;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_157 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_156;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_158 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_157;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_159 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_158;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_160 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_159;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_161 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_160;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_162 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_161;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_163 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_162;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_164 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_163;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_165 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_164;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_166 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_165;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_167 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_166;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_168 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_167;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_169 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_168;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_170 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_169;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_171 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_170;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_172 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_171;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_173 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_172;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_174 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_173;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_175 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_174;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_176 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_175;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_177 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_176;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_178 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_177;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_179 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_178;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_180 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_179;
      dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_181 <= dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98_stage_180;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_138 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_139 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_138;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_140 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_139;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_141 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_140;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_142 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_141;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_143 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_142;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_144 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_143;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_145 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_144;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_146 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_145;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_147 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_146;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_148 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_147;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_149 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_148;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_150 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_149;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_151 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_150;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_152 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_151;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_153 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_152;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_154 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_153;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_155 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_154;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_156 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_155;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_157 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_156;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_158 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_157;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_159 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_158;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_160 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_159;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_161 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_160;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_162 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_161;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_163 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_162;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_164 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_163;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_165 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_164;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_166 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_165;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_167 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_166;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_168 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_167;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_169 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_168;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_170 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_169;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_171 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_170;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_172 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_171;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_173 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_172;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_174 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_173;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_175 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_174;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_176 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_175;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_177 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_176;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_178 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_177;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_179 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_178;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_180 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_179;
      dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_181 <= dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95_stage_180;
      dark_laplace_us_2_update_0_stage_143 <= dark_laplace_us_2_update_0;
      dark_laplace_us_2_update_0_stage_144 <= dark_laplace_us_2_update_0_stage_143;
      dark_laplace_us_2_update_0_stage_145 <= dark_laplace_us_2_update_0_stage_144;
      dark_laplace_us_2_update_0_stage_146 <= dark_laplace_us_2_update_0_stage_145;
      dark_laplace_us_2_update_0_stage_147 <= dark_laplace_us_2_update_0_stage_146;
      dark_laplace_us_2_update_0_stage_148 <= dark_laplace_us_2_update_0_stage_147;
      dark_laplace_us_2_update_0_stage_149 <= dark_laplace_us_2_update_0_stage_148;
      dark_laplace_us_2_update_0_stage_150 <= dark_laplace_us_2_update_0_stage_149;
      dark_laplace_us_2_update_0_stage_151 <= dark_laplace_us_2_update_0_stage_150;
      dark_laplace_us_2_update_0_stage_152 <= dark_laplace_us_2_update_0_stage_151;
      dark_laplace_us_2_update_0_stage_153 <= dark_laplace_us_2_update_0_stage_152;
      dark_laplace_us_2_update_0_stage_154 <= dark_laplace_us_2_update_0_stage_153;
      dark_laplace_us_2_update_0_stage_155 <= dark_laplace_us_2_update_0_stage_154;
      dark_laplace_us_2_update_0_stage_156 <= dark_laplace_us_2_update_0_stage_155;
      dark_laplace_us_2_update_0_stage_157 <= dark_laplace_us_2_update_0_stage_156;
      dark_laplace_us_2_update_0_stage_158 <= dark_laplace_us_2_update_0_stage_157;
      dark_laplace_us_2_update_0_stage_159 <= dark_laplace_us_2_update_0_stage_158;
      dark_laplace_us_2_update_0_stage_160 <= dark_laplace_us_2_update_0_stage_159;
      dark_laplace_us_2_update_0_stage_161 <= dark_laplace_us_2_update_0_stage_160;
      dark_laplace_us_2_update_0_stage_162 <= dark_laplace_us_2_update_0_stage_161;
      dark_laplace_us_2_update_0_stage_163 <= dark_laplace_us_2_update_0_stage_162;
      dark_laplace_us_2_update_0_stage_164 <= dark_laplace_us_2_update_0_stage_163;
      dark_laplace_us_2_update_0_stage_165 <= dark_laplace_us_2_update_0_stage_164;
      dark_laplace_us_2_update_0_stage_166 <= dark_laplace_us_2_update_0_stage_165;
      dark_laplace_us_2_update_0_stage_167 <= dark_laplace_us_2_update_0_stage_166;
      dark_laplace_us_2_update_0_stage_168 <= dark_laplace_us_2_update_0_stage_167;
      dark_laplace_us_2_update_0_stage_169 <= dark_laplace_us_2_update_0_stage_168;
      dark_laplace_us_2_update_0_stage_170 <= dark_laplace_us_2_update_0_stage_169;
      dark_laplace_us_2_update_0_stage_171 <= dark_laplace_us_2_update_0_stage_170;
      dark_laplace_us_2_update_0_stage_172 <= dark_laplace_us_2_update_0_stage_171;
      dark_laplace_us_2_update_0_stage_173 <= dark_laplace_us_2_update_0_stage_172;
      dark_laplace_us_2_update_0_stage_174 <= dark_laplace_us_2_update_0_stage_173;
      dark_laplace_us_2_update_0_stage_175 <= dark_laplace_us_2_update_0_stage_174;
      dark_laplace_us_2_update_0_stage_176 <= dark_laplace_us_2_update_0_stage_175;
      dark_laplace_us_2_update_0_stage_177 <= dark_laplace_us_2_update_0_stage_176;
      dark_laplace_us_2_update_0_stage_178 <= dark_laplace_us_2_update_0_stage_177;
      dark_laplace_us_2_update_0_stage_179 <= dark_laplace_us_2_update_0_stage_178;
      dark_laplace_us_2_update_0_stage_180 <= dark_laplace_us_2_update_0_stage_179;
      dark_laplace_us_2_update_0_stage_181 <= dark_laplace_us_2_update_0_stage_180;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_144 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_145 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_144;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_146 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_145;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_147 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_146;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_148 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_147;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_149 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_148;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_150 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_149;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_151 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_150;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_152 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_151;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_153 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_152;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_154 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_153;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_155 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_154;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_156 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_155;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_157 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_156;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_158 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_157;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_159 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_158;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_160 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_159;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_161 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_160;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_162 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_161;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_163 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_162;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_164 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_163;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_165 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_164;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_166 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_165;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_167 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_166;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_168 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_167;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_169 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_168;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_170 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_169;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_171 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_170;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_172 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_171;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_173 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_172;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_174 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_173;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_175 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_174;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_176 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_175;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_177 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_176;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_178 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_177;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_179 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_178;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_180 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_179;
      dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_181 <= dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99_stage_180;
      final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_179 <= final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126;
      final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_180 <= final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_179;
      final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_181 <= final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126_stage_180;
      pyramid_synthetic_exposure_fusion_update_0_stage_180 <= pyramid_synthetic_exposure_fusion_update_0;
      pyramid_synthetic_exposure_fusion_update_0_stage_181 <= pyramid_synthetic_exposure_fusion_update_0_stage_180;
      pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127_stage_181 <= pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_23 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_24 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_23;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_25 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_24;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_26 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_25;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_27 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_26;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_28 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_27;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_29 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_28;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_30 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_29;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_31 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_30;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_32 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_31;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_33 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_32;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_34 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_33;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_35 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_34;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_36 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_35;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_37 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_36;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_38 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_37;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_39 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_38;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_40 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_39;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_41 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_40;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_42 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_41;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_43 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_42;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_44 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_43;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_45 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_44;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_46 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_45;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_47 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_46;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_48 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_47;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_49 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_48;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_50 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_49;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_51 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_50;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_52 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_51;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_53 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_52;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_54 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_53;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_55 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_54;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_56 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_55;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_57 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_56;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_58 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_57;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_59 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_58;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_60 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_59;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_61 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_60;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_62 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_61;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_63 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_62;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_64 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_63;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_65 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_64;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_66 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_65;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_67 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_66;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_68 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_67;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_69 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_68;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_70 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_69;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_71 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_70;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_72 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_71;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_73 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_72;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_74 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_73;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_75 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_74;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_76 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_75;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_77 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_76;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_78 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_77;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_79 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_78;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_80 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_79;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_81 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_80;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_82 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_81;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_83 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_82;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_84 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_83;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_85 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_84;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_86 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_85;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_87 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_86;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_88 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_87;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_89 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_88;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_90 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_89;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_91 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_90;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_92 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_91;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_93 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_92;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_94 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_93;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_95 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_94;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_96 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_95;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_97 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_96;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_98 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_97;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_99 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_98;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_100 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_99;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_101 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_100;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_102 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_101;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_103 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_102;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_104 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_103;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_105 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_104;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_106 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_105;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_107 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_106;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_108 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_107;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_109 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_108;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_110 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_109;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_111 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_110;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_112 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_111;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_113 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_112;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_114 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_113;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_115 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_114;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_116 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_115;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_117 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_116;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_118 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_117;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_119 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_118;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_120 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_119;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_121 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_120;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_122 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_121;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_123 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_122;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_124 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_123;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_125 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_124;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_126 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_125;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_127 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_126;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_128 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_127;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_129 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_128;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_130 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_129;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_131 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_130;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_132 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_131;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_133 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_132;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_134 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_133;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_135 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_134;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_136 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_135;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_137 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_136;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_138 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_137;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_139 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_138;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_140 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_139;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_141 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_140;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_142 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_141;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_143 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_142;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_144 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_143;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_145 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_144;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_146 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_145;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_147 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_146;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_148 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_147;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_149 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_148;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_150 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_149;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_151 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_150;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_152 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_151;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_153 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_152;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_154 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_153;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_155 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_154;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_156 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_155;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_157 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_156;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_158 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_157;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_159 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_158;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_160 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_159;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_161 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_160;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_162 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_161;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_163 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_162;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_164 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_163;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_165 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_164;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_166 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_165;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_167 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_166;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_168 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_167;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_169 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_168;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_170 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_169;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_171 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_170;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_172 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_171;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_173 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_172;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_174 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_173;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_175 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_174;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_176 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_175;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_177 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_176;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_178 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_177;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_179 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_178;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_180 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_179;
      dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_181 <= dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14_stage_180;
      dark_gauss_ds_1_update_0_stage_24 <= dark_gauss_ds_1_update_0;
      dark_gauss_ds_1_update_0_stage_25 <= dark_gauss_ds_1_update_0_stage_24;
      dark_gauss_ds_1_update_0_stage_26 <= dark_gauss_ds_1_update_0_stage_25;
      dark_gauss_ds_1_update_0_stage_27 <= dark_gauss_ds_1_update_0_stage_26;
      dark_gauss_ds_1_update_0_stage_28 <= dark_gauss_ds_1_update_0_stage_27;
      dark_gauss_ds_1_update_0_stage_29 <= dark_gauss_ds_1_update_0_stage_28;
      dark_gauss_ds_1_update_0_stage_30 <= dark_gauss_ds_1_update_0_stage_29;
      dark_gauss_ds_1_update_0_stage_31 <= dark_gauss_ds_1_update_0_stage_30;
      dark_gauss_ds_1_update_0_stage_32 <= dark_gauss_ds_1_update_0_stage_31;
      dark_gauss_ds_1_update_0_stage_33 <= dark_gauss_ds_1_update_0_stage_32;
      dark_gauss_ds_1_update_0_stage_34 <= dark_gauss_ds_1_update_0_stage_33;
      dark_gauss_ds_1_update_0_stage_35 <= dark_gauss_ds_1_update_0_stage_34;
      dark_gauss_ds_1_update_0_stage_36 <= dark_gauss_ds_1_update_0_stage_35;
      dark_gauss_ds_1_update_0_stage_37 <= dark_gauss_ds_1_update_0_stage_36;
      dark_gauss_ds_1_update_0_stage_38 <= dark_gauss_ds_1_update_0_stage_37;
      dark_gauss_ds_1_update_0_stage_39 <= dark_gauss_ds_1_update_0_stage_38;
      dark_gauss_ds_1_update_0_stage_40 <= dark_gauss_ds_1_update_0_stage_39;
      dark_gauss_ds_1_update_0_stage_41 <= dark_gauss_ds_1_update_0_stage_40;
      dark_gauss_ds_1_update_0_stage_42 <= dark_gauss_ds_1_update_0_stage_41;
      dark_gauss_ds_1_update_0_stage_43 <= dark_gauss_ds_1_update_0_stage_42;
      dark_gauss_ds_1_update_0_stage_44 <= dark_gauss_ds_1_update_0_stage_43;
      dark_gauss_ds_1_update_0_stage_45 <= dark_gauss_ds_1_update_0_stage_44;
      dark_gauss_ds_1_update_0_stage_46 <= dark_gauss_ds_1_update_0_stage_45;
      dark_gauss_ds_1_update_0_stage_47 <= dark_gauss_ds_1_update_0_stage_46;
      dark_gauss_ds_1_update_0_stage_48 <= dark_gauss_ds_1_update_0_stage_47;
      dark_gauss_ds_1_update_0_stage_49 <= dark_gauss_ds_1_update_0_stage_48;
      dark_gauss_ds_1_update_0_stage_50 <= dark_gauss_ds_1_update_0_stage_49;
      dark_gauss_ds_1_update_0_stage_51 <= dark_gauss_ds_1_update_0_stage_50;
      dark_gauss_ds_1_update_0_stage_52 <= dark_gauss_ds_1_update_0_stage_51;
      dark_gauss_ds_1_update_0_stage_53 <= dark_gauss_ds_1_update_0_stage_52;
      dark_gauss_ds_1_update_0_stage_54 <= dark_gauss_ds_1_update_0_stage_53;
      dark_gauss_ds_1_update_0_stage_55 <= dark_gauss_ds_1_update_0_stage_54;
      dark_gauss_ds_1_update_0_stage_56 <= dark_gauss_ds_1_update_0_stage_55;
      dark_gauss_ds_1_update_0_stage_57 <= dark_gauss_ds_1_update_0_stage_56;
      dark_gauss_ds_1_update_0_stage_58 <= dark_gauss_ds_1_update_0_stage_57;
      dark_gauss_ds_1_update_0_stage_59 <= dark_gauss_ds_1_update_0_stage_58;
      dark_gauss_ds_1_update_0_stage_60 <= dark_gauss_ds_1_update_0_stage_59;
      dark_gauss_ds_1_update_0_stage_61 <= dark_gauss_ds_1_update_0_stage_60;
      dark_gauss_ds_1_update_0_stage_62 <= dark_gauss_ds_1_update_0_stage_61;
      dark_gauss_ds_1_update_0_stage_63 <= dark_gauss_ds_1_update_0_stage_62;
      dark_gauss_ds_1_update_0_stage_64 <= dark_gauss_ds_1_update_0_stage_63;
      dark_gauss_ds_1_update_0_stage_65 <= dark_gauss_ds_1_update_0_stage_64;
      dark_gauss_ds_1_update_0_stage_66 <= dark_gauss_ds_1_update_0_stage_65;
      dark_gauss_ds_1_update_0_stage_67 <= dark_gauss_ds_1_update_0_stage_66;
      dark_gauss_ds_1_update_0_stage_68 <= dark_gauss_ds_1_update_0_stage_67;
      dark_gauss_ds_1_update_0_stage_69 <= dark_gauss_ds_1_update_0_stage_68;
      dark_gauss_ds_1_update_0_stage_70 <= dark_gauss_ds_1_update_0_stage_69;
      dark_gauss_ds_1_update_0_stage_71 <= dark_gauss_ds_1_update_0_stage_70;
      dark_gauss_ds_1_update_0_stage_72 <= dark_gauss_ds_1_update_0_stage_71;
      dark_gauss_ds_1_update_0_stage_73 <= dark_gauss_ds_1_update_0_stage_72;
      dark_gauss_ds_1_update_0_stage_74 <= dark_gauss_ds_1_update_0_stage_73;
      dark_gauss_ds_1_update_0_stage_75 <= dark_gauss_ds_1_update_0_stage_74;
      dark_gauss_ds_1_update_0_stage_76 <= dark_gauss_ds_1_update_0_stage_75;
      dark_gauss_ds_1_update_0_stage_77 <= dark_gauss_ds_1_update_0_stage_76;
      dark_gauss_ds_1_update_0_stage_78 <= dark_gauss_ds_1_update_0_stage_77;
      dark_gauss_ds_1_update_0_stage_79 <= dark_gauss_ds_1_update_0_stage_78;
      dark_gauss_ds_1_update_0_stage_80 <= dark_gauss_ds_1_update_0_stage_79;
      dark_gauss_ds_1_update_0_stage_81 <= dark_gauss_ds_1_update_0_stage_80;
      dark_gauss_ds_1_update_0_stage_82 <= dark_gauss_ds_1_update_0_stage_81;
      dark_gauss_ds_1_update_0_stage_83 <= dark_gauss_ds_1_update_0_stage_82;
      dark_gauss_ds_1_update_0_stage_84 <= dark_gauss_ds_1_update_0_stage_83;
      dark_gauss_ds_1_update_0_stage_85 <= dark_gauss_ds_1_update_0_stage_84;
      dark_gauss_ds_1_update_0_stage_86 <= dark_gauss_ds_1_update_0_stage_85;
      dark_gauss_ds_1_update_0_stage_87 <= dark_gauss_ds_1_update_0_stage_86;
      dark_gauss_ds_1_update_0_stage_88 <= dark_gauss_ds_1_update_0_stage_87;
      dark_gauss_ds_1_update_0_stage_89 <= dark_gauss_ds_1_update_0_stage_88;
      dark_gauss_ds_1_update_0_stage_90 <= dark_gauss_ds_1_update_0_stage_89;
      dark_gauss_ds_1_update_0_stage_91 <= dark_gauss_ds_1_update_0_stage_90;
      dark_gauss_ds_1_update_0_stage_92 <= dark_gauss_ds_1_update_0_stage_91;
      dark_gauss_ds_1_update_0_stage_93 <= dark_gauss_ds_1_update_0_stage_92;
      dark_gauss_ds_1_update_0_stage_94 <= dark_gauss_ds_1_update_0_stage_93;
      dark_gauss_ds_1_update_0_stage_95 <= dark_gauss_ds_1_update_0_stage_94;
      dark_gauss_ds_1_update_0_stage_96 <= dark_gauss_ds_1_update_0_stage_95;
      dark_gauss_ds_1_update_0_stage_97 <= dark_gauss_ds_1_update_0_stage_96;
      dark_gauss_ds_1_update_0_stage_98 <= dark_gauss_ds_1_update_0_stage_97;
      dark_gauss_ds_1_update_0_stage_99 <= dark_gauss_ds_1_update_0_stage_98;
      dark_gauss_ds_1_update_0_stage_100 <= dark_gauss_ds_1_update_0_stage_99;
      dark_gauss_ds_1_update_0_stage_101 <= dark_gauss_ds_1_update_0_stage_100;
      dark_gauss_ds_1_update_0_stage_102 <= dark_gauss_ds_1_update_0_stage_101;
      dark_gauss_ds_1_update_0_stage_103 <= dark_gauss_ds_1_update_0_stage_102;
      dark_gauss_ds_1_update_0_stage_104 <= dark_gauss_ds_1_update_0_stage_103;
      dark_gauss_ds_1_update_0_stage_105 <= dark_gauss_ds_1_update_0_stage_104;
      dark_gauss_ds_1_update_0_stage_106 <= dark_gauss_ds_1_update_0_stage_105;
      dark_gauss_ds_1_update_0_stage_107 <= dark_gauss_ds_1_update_0_stage_106;
      dark_gauss_ds_1_update_0_stage_108 <= dark_gauss_ds_1_update_0_stage_107;
      dark_gauss_ds_1_update_0_stage_109 <= dark_gauss_ds_1_update_0_stage_108;
      dark_gauss_ds_1_update_0_stage_110 <= dark_gauss_ds_1_update_0_stage_109;
      dark_gauss_ds_1_update_0_stage_111 <= dark_gauss_ds_1_update_0_stage_110;
      dark_gauss_ds_1_update_0_stage_112 <= dark_gauss_ds_1_update_0_stage_111;
      dark_gauss_ds_1_update_0_stage_113 <= dark_gauss_ds_1_update_0_stage_112;
      dark_gauss_ds_1_update_0_stage_114 <= dark_gauss_ds_1_update_0_stage_113;
      dark_gauss_ds_1_update_0_stage_115 <= dark_gauss_ds_1_update_0_stage_114;
      dark_gauss_ds_1_update_0_stage_116 <= dark_gauss_ds_1_update_0_stage_115;
      dark_gauss_ds_1_update_0_stage_117 <= dark_gauss_ds_1_update_0_stage_116;
      dark_gauss_ds_1_update_0_stage_118 <= dark_gauss_ds_1_update_0_stage_117;
      dark_gauss_ds_1_update_0_stage_119 <= dark_gauss_ds_1_update_0_stage_118;
      dark_gauss_ds_1_update_0_stage_120 <= dark_gauss_ds_1_update_0_stage_119;
      dark_gauss_ds_1_update_0_stage_121 <= dark_gauss_ds_1_update_0_stage_120;
      dark_gauss_ds_1_update_0_stage_122 <= dark_gauss_ds_1_update_0_stage_121;
      dark_gauss_ds_1_update_0_stage_123 <= dark_gauss_ds_1_update_0_stage_122;
      dark_gauss_ds_1_update_0_stage_124 <= dark_gauss_ds_1_update_0_stage_123;
      dark_gauss_ds_1_update_0_stage_125 <= dark_gauss_ds_1_update_0_stage_124;
      dark_gauss_ds_1_update_0_stage_126 <= dark_gauss_ds_1_update_0_stage_125;
      dark_gauss_ds_1_update_0_stage_127 <= dark_gauss_ds_1_update_0_stage_126;
      dark_gauss_ds_1_update_0_stage_128 <= dark_gauss_ds_1_update_0_stage_127;
      dark_gauss_ds_1_update_0_stage_129 <= dark_gauss_ds_1_update_0_stage_128;
      dark_gauss_ds_1_update_0_stage_130 <= dark_gauss_ds_1_update_0_stage_129;
      dark_gauss_ds_1_update_0_stage_131 <= dark_gauss_ds_1_update_0_stage_130;
      dark_gauss_ds_1_update_0_stage_132 <= dark_gauss_ds_1_update_0_stage_131;
      dark_gauss_ds_1_update_0_stage_133 <= dark_gauss_ds_1_update_0_stage_132;
      dark_gauss_ds_1_update_0_stage_134 <= dark_gauss_ds_1_update_0_stage_133;
      dark_gauss_ds_1_update_0_stage_135 <= dark_gauss_ds_1_update_0_stage_134;
      dark_gauss_ds_1_update_0_stage_136 <= dark_gauss_ds_1_update_0_stage_135;
      dark_gauss_ds_1_update_0_stage_137 <= dark_gauss_ds_1_update_0_stage_136;
      dark_gauss_ds_1_update_0_stage_138 <= dark_gauss_ds_1_update_0_stage_137;
      dark_gauss_ds_1_update_0_stage_139 <= dark_gauss_ds_1_update_0_stage_138;
      dark_gauss_ds_1_update_0_stage_140 <= dark_gauss_ds_1_update_0_stage_139;
      dark_gauss_ds_1_update_0_stage_141 <= dark_gauss_ds_1_update_0_stage_140;
      dark_gauss_ds_1_update_0_stage_142 <= dark_gauss_ds_1_update_0_stage_141;
      dark_gauss_ds_1_update_0_stage_143 <= dark_gauss_ds_1_update_0_stage_142;
      dark_gauss_ds_1_update_0_stage_144 <= dark_gauss_ds_1_update_0_stage_143;
      dark_gauss_ds_1_update_0_stage_145 <= dark_gauss_ds_1_update_0_stage_144;
      dark_gauss_ds_1_update_0_stage_146 <= dark_gauss_ds_1_update_0_stage_145;
      dark_gauss_ds_1_update_0_stage_147 <= dark_gauss_ds_1_update_0_stage_146;
      dark_gauss_ds_1_update_0_stage_148 <= dark_gauss_ds_1_update_0_stage_147;
      dark_gauss_ds_1_update_0_stage_149 <= dark_gauss_ds_1_update_0_stage_148;
      dark_gauss_ds_1_update_0_stage_150 <= dark_gauss_ds_1_update_0_stage_149;
      dark_gauss_ds_1_update_0_stage_151 <= dark_gauss_ds_1_update_0_stage_150;
      dark_gauss_ds_1_update_0_stage_152 <= dark_gauss_ds_1_update_0_stage_151;
      dark_gauss_ds_1_update_0_stage_153 <= dark_gauss_ds_1_update_0_stage_152;
      dark_gauss_ds_1_update_0_stage_154 <= dark_gauss_ds_1_update_0_stage_153;
      dark_gauss_ds_1_update_0_stage_155 <= dark_gauss_ds_1_update_0_stage_154;
      dark_gauss_ds_1_update_0_stage_156 <= dark_gauss_ds_1_update_0_stage_155;
      dark_gauss_ds_1_update_0_stage_157 <= dark_gauss_ds_1_update_0_stage_156;
      dark_gauss_ds_1_update_0_stage_158 <= dark_gauss_ds_1_update_0_stage_157;
      dark_gauss_ds_1_update_0_stage_159 <= dark_gauss_ds_1_update_0_stage_158;
      dark_gauss_ds_1_update_0_stage_160 <= dark_gauss_ds_1_update_0_stage_159;
      dark_gauss_ds_1_update_0_stage_161 <= dark_gauss_ds_1_update_0_stage_160;
      dark_gauss_ds_1_update_0_stage_162 <= dark_gauss_ds_1_update_0_stage_161;
      dark_gauss_ds_1_update_0_stage_163 <= dark_gauss_ds_1_update_0_stage_162;
      dark_gauss_ds_1_update_0_stage_164 <= dark_gauss_ds_1_update_0_stage_163;
      dark_gauss_ds_1_update_0_stage_165 <= dark_gauss_ds_1_update_0_stage_164;
      dark_gauss_ds_1_update_0_stage_166 <= dark_gauss_ds_1_update_0_stage_165;
      dark_gauss_ds_1_update_0_stage_167 <= dark_gauss_ds_1_update_0_stage_166;
      dark_gauss_ds_1_update_0_stage_168 <= dark_gauss_ds_1_update_0_stage_167;
      dark_gauss_ds_1_update_0_stage_169 <= dark_gauss_ds_1_update_0_stage_168;
      dark_gauss_ds_1_update_0_stage_170 <= dark_gauss_ds_1_update_0_stage_169;
      dark_gauss_ds_1_update_0_stage_171 <= dark_gauss_ds_1_update_0_stage_170;
      dark_gauss_ds_1_update_0_stage_172 <= dark_gauss_ds_1_update_0_stage_171;
      dark_gauss_ds_1_update_0_stage_173 <= dark_gauss_ds_1_update_0_stage_172;
      dark_gauss_ds_1_update_0_stage_174 <= dark_gauss_ds_1_update_0_stage_173;
      dark_gauss_ds_1_update_0_stage_175 <= dark_gauss_ds_1_update_0_stage_174;
      dark_gauss_ds_1_update_0_stage_176 <= dark_gauss_ds_1_update_0_stage_175;
      dark_gauss_ds_1_update_0_stage_177 <= dark_gauss_ds_1_update_0_stage_176;
      dark_gauss_ds_1_update_0_stage_178 <= dark_gauss_ds_1_update_0_stage_177;
      dark_gauss_ds_1_update_0_stage_179 <= dark_gauss_ds_1_update_0_stage_178;
      dark_gauss_ds_1_update_0_stage_180 <= dark_gauss_ds_1_update_0_stage_179;
      dark_gauss_ds_1_update_0_stage_181 <= dark_gauss_ds_1_update_0_stage_180;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_25 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_26 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_25;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_27 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_26;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_28 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_27;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_29 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_28;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_30 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_29;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_31 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_30;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_32 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_31;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_33 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_32;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_34 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_33;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_35 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_34;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_36 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_35;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_37 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_36;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_38 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_37;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_39 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_38;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_40 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_39;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_41 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_40;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_42 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_41;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_43 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_42;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_44 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_43;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_45 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_44;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_46 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_45;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_47 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_46;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_48 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_47;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_49 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_48;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_50 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_49;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_51 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_50;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_52 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_51;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_53 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_52;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_54 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_53;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_55 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_54;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_56 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_55;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_57 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_56;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_58 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_57;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_59 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_58;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_60 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_59;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_61 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_60;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_62 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_61;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_63 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_62;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_64 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_63;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_65 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_64;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_66 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_65;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_67 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_66;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_68 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_67;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_69 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_68;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_70 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_69;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_71 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_70;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_72 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_71;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_73 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_72;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_74 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_73;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_75 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_74;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_76 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_75;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_77 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_76;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_78 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_77;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_79 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_78;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_80 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_79;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_81 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_80;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_82 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_81;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_83 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_82;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_84 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_83;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_85 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_84;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_86 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_85;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_87 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_86;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_88 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_87;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_89 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_88;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_90 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_89;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_91 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_90;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_92 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_91;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_93 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_92;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_94 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_93;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_95 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_94;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_96 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_95;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_97 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_96;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_98 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_97;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_99 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_98;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_100 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_99;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_101 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_100;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_102 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_101;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_103 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_102;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_104 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_103;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_105 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_104;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_106 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_105;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_107 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_106;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_108 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_107;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_109 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_108;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_110 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_109;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_111 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_110;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_112 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_111;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_113 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_112;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_114 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_113;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_115 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_114;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_116 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_115;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_117 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_116;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_118 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_117;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_119 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_118;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_120 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_119;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_121 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_120;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_122 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_121;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_123 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_122;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_124 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_123;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_125 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_124;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_126 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_125;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_127 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_126;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_128 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_127;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_129 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_128;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_130 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_129;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_131 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_130;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_132 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_131;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_133 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_132;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_134 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_133;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_135 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_134;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_136 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_135;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_137 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_136;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_138 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_137;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_139 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_138;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_140 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_139;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_141 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_140;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_142 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_141;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_143 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_142;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_144 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_143;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_145 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_144;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_146 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_145;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_147 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_146;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_148 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_147;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_149 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_148;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_150 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_149;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_151 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_150;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_152 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_151;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_153 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_152;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_154 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_153;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_155 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_154;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_156 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_155;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_157 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_156;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_158 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_157;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_159 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_158;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_160 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_159;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_161 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_160;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_162 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_161;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_163 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_162;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_164 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_163;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_165 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_164;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_166 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_165;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_167 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_166;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_168 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_167;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_169 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_168;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_170 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_169;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_171 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_170;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_172 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_171;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_173 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_172;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_174 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_173;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_175 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_174;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_176 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_175;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_177 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_176;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_178 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_177;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_179 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_178;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_180 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_179;
      dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_181 <= dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15_stage_180;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_31 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_32 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_31;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_33 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_32;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_34 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_33;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_35 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_34;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_36 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_35;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_37 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_36;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_38 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_37;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_39 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_38;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_40 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_39;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_41 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_40;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_42 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_41;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_43 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_42;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_44 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_43;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_45 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_44;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_46 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_45;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_47 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_46;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_48 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_47;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_49 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_48;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_50 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_49;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_51 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_50;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_52 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_51;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_53 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_52;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_54 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_53;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_55 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_54;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_56 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_55;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_57 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_56;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_58 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_57;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_59 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_58;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_60 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_59;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_61 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_60;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_62 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_61;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_63 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_62;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_64 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_63;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_65 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_64;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_66 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_65;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_67 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_66;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_68 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_67;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_69 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_68;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_70 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_69;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_71 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_70;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_72 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_71;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_73 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_72;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_74 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_73;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_75 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_74;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_76 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_75;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_77 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_76;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_78 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_77;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_79 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_78;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_80 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_79;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_81 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_80;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_82 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_81;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_83 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_82;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_84 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_83;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_85 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_84;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_86 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_85;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_87 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_86;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_88 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_87;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_89 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_88;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_90 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_89;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_91 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_90;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_92 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_91;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_93 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_92;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_94 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_93;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_95 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_94;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_96 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_95;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_97 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_96;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_98 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_97;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_99 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_98;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_100 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_99;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_101 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_100;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_102 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_101;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_103 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_102;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_104 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_103;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_105 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_104;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_106 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_105;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_107 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_106;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_108 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_107;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_109 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_108;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_110 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_109;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_111 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_110;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_112 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_111;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_113 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_112;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_114 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_113;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_115 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_114;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_116 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_115;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_117 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_116;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_118 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_117;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_119 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_118;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_120 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_119;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_121 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_120;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_122 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_121;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_123 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_122;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_124 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_123;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_125 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_124;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_126 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_125;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_127 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_126;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_128 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_127;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_129 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_128;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_130 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_129;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_131 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_130;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_132 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_131;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_133 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_132;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_134 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_133;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_135 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_134;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_136 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_135;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_137 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_136;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_138 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_137;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_139 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_138;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_140 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_139;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_141 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_140;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_142 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_141;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_143 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_142;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_144 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_143;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_145 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_144;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_146 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_145;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_147 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_146;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_148 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_147;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_149 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_148;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_150 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_149;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_151 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_150;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_152 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_151;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_153 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_152;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_154 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_153;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_155 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_154;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_156 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_155;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_157 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_156;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_158 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_157;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_159 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_158;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_160 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_159;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_161 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_160;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_162 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_161;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_163 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_162;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_164 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_163;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_165 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_164;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_166 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_165;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_167 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_166;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_168 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_167;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_169 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_168;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_170 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_169;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_171 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_170;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_172 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_171;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_173 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_172;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_174 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_173;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_175 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_174;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_176 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_175;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_177 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_176;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_178 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_177;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_179 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_178;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_180 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_179;
      dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_181 <= dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19_stage_180;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_32 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_33 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_32;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_34 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_33;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_35 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_34;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_36 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_35;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_37 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_36;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_38 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_37;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_39 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_38;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_40 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_39;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_41 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_40;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_42 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_41;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_43 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_42;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_44 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_43;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_45 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_44;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_46 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_45;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_47 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_46;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_48 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_47;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_49 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_48;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_50 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_49;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_51 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_50;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_52 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_51;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_53 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_52;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_54 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_53;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_55 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_54;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_56 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_55;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_57 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_56;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_58 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_57;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_59 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_58;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_60 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_59;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_61 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_60;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_62 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_61;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_63 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_62;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_64 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_63;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_65 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_64;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_66 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_65;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_67 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_66;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_68 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_67;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_69 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_68;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_70 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_69;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_71 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_70;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_72 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_71;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_73 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_72;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_74 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_73;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_75 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_74;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_76 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_75;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_77 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_76;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_78 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_77;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_79 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_78;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_80 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_79;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_81 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_80;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_82 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_81;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_83 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_82;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_84 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_83;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_85 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_84;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_86 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_85;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_87 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_86;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_88 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_87;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_89 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_88;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_90 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_89;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_91 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_90;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_92 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_91;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_93 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_92;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_94 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_93;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_95 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_94;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_96 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_95;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_97 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_96;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_98 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_97;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_99 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_98;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_100 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_99;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_101 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_100;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_102 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_101;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_103 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_102;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_104 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_103;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_105 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_104;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_106 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_105;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_107 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_106;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_108 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_107;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_109 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_108;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_110 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_109;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_111 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_110;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_112 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_111;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_113 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_112;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_114 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_113;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_115 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_114;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_116 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_115;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_117 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_116;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_118 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_117;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_119 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_118;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_120 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_119;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_121 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_120;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_122 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_121;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_123 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_122;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_124 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_123;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_125 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_124;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_126 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_125;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_127 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_126;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_128 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_127;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_129 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_128;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_130 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_129;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_131 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_130;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_132 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_131;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_133 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_132;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_134 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_133;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_135 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_134;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_136 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_135;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_137 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_136;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_138 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_137;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_139 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_138;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_140 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_139;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_141 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_140;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_142 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_141;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_143 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_142;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_144 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_143;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_145 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_144;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_146 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_145;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_147 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_146;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_148 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_147;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_149 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_148;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_150 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_149;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_151 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_150;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_152 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_151;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_153 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_152;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_154 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_153;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_155 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_154;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_156 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_155;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_157 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_156;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_158 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_157;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_159 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_158;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_160 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_159;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_161 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_160;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_162 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_161;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_163 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_162;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_164 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_163;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_165 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_164;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_166 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_165;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_167 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_166;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_168 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_167;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_169 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_168;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_170 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_169;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_171 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_170;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_172 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_171;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_173 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_172;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_174 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_173;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_175 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_174;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_176 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_175;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_177 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_176;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_178 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_177;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_179 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_178;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_180 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_179;
      bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_181 <= bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20_stage_180;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_29 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_30 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_29;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_31 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_30;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_32 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_31;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_33 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_32;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_34 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_33;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_35 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_34;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_36 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_35;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_37 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_36;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_38 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_37;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_39 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_38;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_40 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_39;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_41 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_40;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_42 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_41;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_43 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_42;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_44 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_43;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_45 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_44;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_46 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_45;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_47 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_46;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_48 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_47;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_49 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_48;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_50 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_49;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_51 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_50;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_52 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_51;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_53 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_52;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_54 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_53;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_55 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_54;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_56 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_55;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_57 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_56;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_58 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_57;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_59 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_58;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_60 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_59;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_61 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_60;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_62 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_61;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_63 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_62;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_64 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_63;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_65 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_64;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_66 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_65;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_67 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_66;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_68 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_67;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_69 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_68;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_70 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_69;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_71 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_70;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_72 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_71;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_73 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_72;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_74 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_73;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_75 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_74;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_76 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_75;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_77 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_76;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_78 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_77;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_79 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_78;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_80 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_79;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_81 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_80;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_82 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_81;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_83 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_82;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_84 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_83;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_85 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_84;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_86 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_85;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_87 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_86;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_88 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_87;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_89 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_88;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_90 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_89;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_91 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_90;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_92 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_91;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_93 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_92;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_94 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_93;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_95 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_94;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_96 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_95;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_97 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_96;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_98 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_97;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_99 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_98;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_100 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_99;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_101 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_100;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_102 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_101;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_103 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_102;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_104 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_103;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_105 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_104;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_106 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_105;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_107 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_106;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_108 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_107;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_109 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_108;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_110 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_109;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_111 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_110;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_112 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_111;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_113 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_112;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_114 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_113;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_115 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_114;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_116 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_115;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_117 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_116;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_118 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_117;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_119 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_118;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_120 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_119;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_121 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_120;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_122 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_121;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_123 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_122;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_124 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_123;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_125 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_124;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_126 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_125;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_127 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_126;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_128 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_127;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_129 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_128;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_130 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_129;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_131 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_130;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_132 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_131;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_133 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_132;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_134 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_133;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_135 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_134;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_136 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_135;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_137 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_136;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_138 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_137;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_139 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_138;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_140 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_139;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_141 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_140;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_142 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_141;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_143 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_142;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_144 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_143;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_145 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_144;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_146 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_145;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_147 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_146;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_148 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_147;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_149 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_148;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_150 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_149;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_151 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_150;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_152 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_151;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_153 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_152;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_154 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_153;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_155 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_154;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_156 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_155;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_157 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_156;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_158 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_157;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_159 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_158;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_160 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_159;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_161 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_160;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_162 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_161;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_163 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_162;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_164 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_163;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_165 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_164;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_166 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_165;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_167 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_166;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_168 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_167;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_169 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_168;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_170 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_169;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_171 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_170;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_172 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_171;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_173 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_172;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_174 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_173;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_175 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_174;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_176 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_175;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_177 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_176;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_178 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_177;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_179 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_178;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_180 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_179;
      dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_181 <= dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18_stage_180;
      dark_gauss_blur_2_update_0_stage_30 <= dark_gauss_blur_2_update_0;
      dark_gauss_blur_2_update_0_stage_31 <= dark_gauss_blur_2_update_0_stage_30;
      dark_gauss_blur_2_update_0_stage_32 <= dark_gauss_blur_2_update_0_stage_31;
      dark_gauss_blur_2_update_0_stage_33 <= dark_gauss_blur_2_update_0_stage_32;
      dark_gauss_blur_2_update_0_stage_34 <= dark_gauss_blur_2_update_0_stage_33;
      dark_gauss_blur_2_update_0_stage_35 <= dark_gauss_blur_2_update_0_stage_34;
      dark_gauss_blur_2_update_0_stage_36 <= dark_gauss_blur_2_update_0_stage_35;
      dark_gauss_blur_2_update_0_stage_37 <= dark_gauss_blur_2_update_0_stage_36;
      dark_gauss_blur_2_update_0_stage_38 <= dark_gauss_blur_2_update_0_stage_37;
      dark_gauss_blur_2_update_0_stage_39 <= dark_gauss_blur_2_update_0_stage_38;
      dark_gauss_blur_2_update_0_stage_40 <= dark_gauss_blur_2_update_0_stage_39;
      dark_gauss_blur_2_update_0_stage_41 <= dark_gauss_blur_2_update_0_stage_40;
      dark_gauss_blur_2_update_0_stage_42 <= dark_gauss_blur_2_update_0_stage_41;
      dark_gauss_blur_2_update_0_stage_43 <= dark_gauss_blur_2_update_0_stage_42;
      dark_gauss_blur_2_update_0_stage_44 <= dark_gauss_blur_2_update_0_stage_43;
      dark_gauss_blur_2_update_0_stage_45 <= dark_gauss_blur_2_update_0_stage_44;
      dark_gauss_blur_2_update_0_stage_46 <= dark_gauss_blur_2_update_0_stage_45;
      dark_gauss_blur_2_update_0_stage_47 <= dark_gauss_blur_2_update_0_stage_46;
      dark_gauss_blur_2_update_0_stage_48 <= dark_gauss_blur_2_update_0_stage_47;
      dark_gauss_blur_2_update_0_stage_49 <= dark_gauss_blur_2_update_0_stage_48;
      dark_gauss_blur_2_update_0_stage_50 <= dark_gauss_blur_2_update_0_stage_49;
      dark_gauss_blur_2_update_0_stage_51 <= dark_gauss_blur_2_update_0_stage_50;
      dark_gauss_blur_2_update_0_stage_52 <= dark_gauss_blur_2_update_0_stage_51;
      dark_gauss_blur_2_update_0_stage_53 <= dark_gauss_blur_2_update_0_stage_52;
      dark_gauss_blur_2_update_0_stage_54 <= dark_gauss_blur_2_update_0_stage_53;
      dark_gauss_blur_2_update_0_stage_55 <= dark_gauss_blur_2_update_0_stage_54;
      dark_gauss_blur_2_update_0_stage_56 <= dark_gauss_blur_2_update_0_stage_55;
      dark_gauss_blur_2_update_0_stage_57 <= dark_gauss_blur_2_update_0_stage_56;
      dark_gauss_blur_2_update_0_stage_58 <= dark_gauss_blur_2_update_0_stage_57;
      dark_gauss_blur_2_update_0_stage_59 <= dark_gauss_blur_2_update_0_stage_58;
      dark_gauss_blur_2_update_0_stage_60 <= dark_gauss_blur_2_update_0_stage_59;
      dark_gauss_blur_2_update_0_stage_61 <= dark_gauss_blur_2_update_0_stage_60;
      dark_gauss_blur_2_update_0_stage_62 <= dark_gauss_blur_2_update_0_stage_61;
      dark_gauss_blur_2_update_0_stage_63 <= dark_gauss_blur_2_update_0_stage_62;
      dark_gauss_blur_2_update_0_stage_64 <= dark_gauss_blur_2_update_0_stage_63;
      dark_gauss_blur_2_update_0_stage_65 <= dark_gauss_blur_2_update_0_stage_64;
      dark_gauss_blur_2_update_0_stage_66 <= dark_gauss_blur_2_update_0_stage_65;
      dark_gauss_blur_2_update_0_stage_67 <= dark_gauss_blur_2_update_0_stage_66;
      dark_gauss_blur_2_update_0_stage_68 <= dark_gauss_blur_2_update_0_stage_67;
      dark_gauss_blur_2_update_0_stage_69 <= dark_gauss_blur_2_update_0_stage_68;
      dark_gauss_blur_2_update_0_stage_70 <= dark_gauss_blur_2_update_0_stage_69;
      dark_gauss_blur_2_update_0_stage_71 <= dark_gauss_blur_2_update_0_stage_70;
      dark_gauss_blur_2_update_0_stage_72 <= dark_gauss_blur_2_update_0_stage_71;
      dark_gauss_blur_2_update_0_stage_73 <= dark_gauss_blur_2_update_0_stage_72;
      dark_gauss_blur_2_update_0_stage_74 <= dark_gauss_blur_2_update_0_stage_73;
      dark_gauss_blur_2_update_0_stage_75 <= dark_gauss_blur_2_update_0_stage_74;
      dark_gauss_blur_2_update_0_stage_76 <= dark_gauss_blur_2_update_0_stage_75;
      dark_gauss_blur_2_update_0_stage_77 <= dark_gauss_blur_2_update_0_stage_76;
      dark_gauss_blur_2_update_0_stage_78 <= dark_gauss_blur_2_update_0_stage_77;
      dark_gauss_blur_2_update_0_stage_79 <= dark_gauss_blur_2_update_0_stage_78;
      dark_gauss_blur_2_update_0_stage_80 <= dark_gauss_blur_2_update_0_stage_79;
      dark_gauss_blur_2_update_0_stage_81 <= dark_gauss_blur_2_update_0_stage_80;
      dark_gauss_blur_2_update_0_stage_82 <= dark_gauss_blur_2_update_0_stage_81;
      dark_gauss_blur_2_update_0_stage_83 <= dark_gauss_blur_2_update_0_stage_82;
      dark_gauss_blur_2_update_0_stage_84 <= dark_gauss_blur_2_update_0_stage_83;
      dark_gauss_blur_2_update_0_stage_85 <= dark_gauss_blur_2_update_0_stage_84;
      dark_gauss_blur_2_update_0_stage_86 <= dark_gauss_blur_2_update_0_stage_85;
      dark_gauss_blur_2_update_0_stage_87 <= dark_gauss_blur_2_update_0_stage_86;
      dark_gauss_blur_2_update_0_stage_88 <= dark_gauss_blur_2_update_0_stage_87;
      dark_gauss_blur_2_update_0_stage_89 <= dark_gauss_blur_2_update_0_stage_88;
      dark_gauss_blur_2_update_0_stage_90 <= dark_gauss_blur_2_update_0_stage_89;
      dark_gauss_blur_2_update_0_stage_91 <= dark_gauss_blur_2_update_0_stage_90;
      dark_gauss_blur_2_update_0_stage_92 <= dark_gauss_blur_2_update_0_stage_91;
      dark_gauss_blur_2_update_0_stage_93 <= dark_gauss_blur_2_update_0_stage_92;
      dark_gauss_blur_2_update_0_stage_94 <= dark_gauss_blur_2_update_0_stage_93;
      dark_gauss_blur_2_update_0_stage_95 <= dark_gauss_blur_2_update_0_stage_94;
      dark_gauss_blur_2_update_0_stage_96 <= dark_gauss_blur_2_update_0_stage_95;
      dark_gauss_blur_2_update_0_stage_97 <= dark_gauss_blur_2_update_0_stage_96;
      dark_gauss_blur_2_update_0_stage_98 <= dark_gauss_blur_2_update_0_stage_97;
      dark_gauss_blur_2_update_0_stage_99 <= dark_gauss_blur_2_update_0_stage_98;
      dark_gauss_blur_2_update_0_stage_100 <= dark_gauss_blur_2_update_0_stage_99;
      dark_gauss_blur_2_update_0_stage_101 <= dark_gauss_blur_2_update_0_stage_100;
      dark_gauss_blur_2_update_0_stage_102 <= dark_gauss_blur_2_update_0_stage_101;
      dark_gauss_blur_2_update_0_stage_103 <= dark_gauss_blur_2_update_0_stage_102;
      dark_gauss_blur_2_update_0_stage_104 <= dark_gauss_blur_2_update_0_stage_103;
      dark_gauss_blur_2_update_0_stage_105 <= dark_gauss_blur_2_update_0_stage_104;
      dark_gauss_blur_2_update_0_stage_106 <= dark_gauss_blur_2_update_0_stage_105;
      dark_gauss_blur_2_update_0_stage_107 <= dark_gauss_blur_2_update_0_stage_106;
      dark_gauss_blur_2_update_0_stage_108 <= dark_gauss_blur_2_update_0_stage_107;
      dark_gauss_blur_2_update_0_stage_109 <= dark_gauss_blur_2_update_0_stage_108;
      dark_gauss_blur_2_update_0_stage_110 <= dark_gauss_blur_2_update_0_stage_109;
      dark_gauss_blur_2_update_0_stage_111 <= dark_gauss_blur_2_update_0_stage_110;
      dark_gauss_blur_2_update_0_stage_112 <= dark_gauss_blur_2_update_0_stage_111;
      dark_gauss_blur_2_update_0_stage_113 <= dark_gauss_blur_2_update_0_stage_112;
      dark_gauss_blur_2_update_0_stage_114 <= dark_gauss_blur_2_update_0_stage_113;
      dark_gauss_blur_2_update_0_stage_115 <= dark_gauss_blur_2_update_0_stage_114;
      dark_gauss_blur_2_update_0_stage_116 <= dark_gauss_blur_2_update_0_stage_115;
      dark_gauss_blur_2_update_0_stage_117 <= dark_gauss_blur_2_update_0_stage_116;
      dark_gauss_blur_2_update_0_stage_118 <= dark_gauss_blur_2_update_0_stage_117;
      dark_gauss_blur_2_update_0_stage_119 <= dark_gauss_blur_2_update_0_stage_118;
      dark_gauss_blur_2_update_0_stage_120 <= dark_gauss_blur_2_update_0_stage_119;
      dark_gauss_blur_2_update_0_stage_121 <= dark_gauss_blur_2_update_0_stage_120;
      dark_gauss_blur_2_update_0_stage_122 <= dark_gauss_blur_2_update_0_stage_121;
      dark_gauss_blur_2_update_0_stage_123 <= dark_gauss_blur_2_update_0_stage_122;
      dark_gauss_blur_2_update_0_stage_124 <= dark_gauss_blur_2_update_0_stage_123;
      dark_gauss_blur_2_update_0_stage_125 <= dark_gauss_blur_2_update_0_stage_124;
      dark_gauss_blur_2_update_0_stage_126 <= dark_gauss_blur_2_update_0_stage_125;
      dark_gauss_blur_2_update_0_stage_127 <= dark_gauss_blur_2_update_0_stage_126;
      dark_gauss_blur_2_update_0_stage_128 <= dark_gauss_blur_2_update_0_stage_127;
      dark_gauss_blur_2_update_0_stage_129 <= dark_gauss_blur_2_update_0_stage_128;
      dark_gauss_blur_2_update_0_stage_130 <= dark_gauss_blur_2_update_0_stage_129;
      dark_gauss_blur_2_update_0_stage_131 <= dark_gauss_blur_2_update_0_stage_130;
      dark_gauss_blur_2_update_0_stage_132 <= dark_gauss_blur_2_update_0_stage_131;
      dark_gauss_blur_2_update_0_stage_133 <= dark_gauss_blur_2_update_0_stage_132;
      dark_gauss_blur_2_update_0_stage_134 <= dark_gauss_blur_2_update_0_stage_133;
      dark_gauss_blur_2_update_0_stage_135 <= dark_gauss_blur_2_update_0_stage_134;
      dark_gauss_blur_2_update_0_stage_136 <= dark_gauss_blur_2_update_0_stage_135;
      dark_gauss_blur_2_update_0_stage_137 <= dark_gauss_blur_2_update_0_stage_136;
      dark_gauss_blur_2_update_0_stage_138 <= dark_gauss_blur_2_update_0_stage_137;
      dark_gauss_blur_2_update_0_stage_139 <= dark_gauss_blur_2_update_0_stage_138;
      dark_gauss_blur_2_update_0_stage_140 <= dark_gauss_blur_2_update_0_stage_139;
      dark_gauss_blur_2_update_0_stage_141 <= dark_gauss_blur_2_update_0_stage_140;
      dark_gauss_blur_2_update_0_stage_142 <= dark_gauss_blur_2_update_0_stage_141;
      dark_gauss_blur_2_update_0_stage_143 <= dark_gauss_blur_2_update_0_stage_142;
      dark_gauss_blur_2_update_0_stage_144 <= dark_gauss_blur_2_update_0_stage_143;
      dark_gauss_blur_2_update_0_stage_145 <= dark_gauss_blur_2_update_0_stage_144;
      dark_gauss_blur_2_update_0_stage_146 <= dark_gauss_blur_2_update_0_stage_145;
      dark_gauss_blur_2_update_0_stage_147 <= dark_gauss_blur_2_update_0_stage_146;
      dark_gauss_blur_2_update_0_stage_148 <= dark_gauss_blur_2_update_0_stage_147;
      dark_gauss_blur_2_update_0_stage_149 <= dark_gauss_blur_2_update_0_stage_148;
      dark_gauss_blur_2_update_0_stage_150 <= dark_gauss_blur_2_update_0_stage_149;
      dark_gauss_blur_2_update_0_stage_151 <= dark_gauss_blur_2_update_0_stage_150;
      dark_gauss_blur_2_update_0_stage_152 <= dark_gauss_blur_2_update_0_stage_151;
      dark_gauss_blur_2_update_0_stage_153 <= dark_gauss_blur_2_update_0_stage_152;
      dark_gauss_blur_2_update_0_stage_154 <= dark_gauss_blur_2_update_0_stage_153;
      dark_gauss_blur_2_update_0_stage_155 <= dark_gauss_blur_2_update_0_stage_154;
      dark_gauss_blur_2_update_0_stage_156 <= dark_gauss_blur_2_update_0_stage_155;
      dark_gauss_blur_2_update_0_stage_157 <= dark_gauss_blur_2_update_0_stage_156;
      dark_gauss_blur_2_update_0_stage_158 <= dark_gauss_blur_2_update_0_stage_157;
      dark_gauss_blur_2_update_0_stage_159 <= dark_gauss_blur_2_update_0_stage_158;
      dark_gauss_blur_2_update_0_stage_160 <= dark_gauss_blur_2_update_0_stage_159;
      dark_gauss_blur_2_update_0_stage_161 <= dark_gauss_blur_2_update_0_stage_160;
      dark_gauss_blur_2_update_0_stage_162 <= dark_gauss_blur_2_update_0_stage_161;
      dark_gauss_blur_2_update_0_stage_163 <= dark_gauss_blur_2_update_0_stage_162;
      dark_gauss_blur_2_update_0_stage_164 <= dark_gauss_blur_2_update_0_stage_163;
      dark_gauss_blur_2_update_0_stage_165 <= dark_gauss_blur_2_update_0_stage_164;
      dark_gauss_blur_2_update_0_stage_166 <= dark_gauss_blur_2_update_0_stage_165;
      dark_gauss_blur_2_update_0_stage_167 <= dark_gauss_blur_2_update_0_stage_166;
      dark_gauss_blur_2_update_0_stage_168 <= dark_gauss_blur_2_update_0_stage_167;
      dark_gauss_blur_2_update_0_stage_169 <= dark_gauss_blur_2_update_0_stage_168;
      dark_gauss_blur_2_update_0_stage_170 <= dark_gauss_blur_2_update_0_stage_169;
      dark_gauss_blur_2_update_0_stage_171 <= dark_gauss_blur_2_update_0_stage_170;
      dark_gauss_blur_2_update_0_stage_172 <= dark_gauss_blur_2_update_0_stage_171;
      dark_gauss_blur_2_update_0_stage_173 <= dark_gauss_blur_2_update_0_stage_172;
      dark_gauss_blur_2_update_0_stage_174 <= dark_gauss_blur_2_update_0_stage_173;
      dark_gauss_blur_2_update_0_stage_175 <= dark_gauss_blur_2_update_0_stage_174;
      dark_gauss_blur_2_update_0_stage_176 <= dark_gauss_blur_2_update_0_stage_175;
      dark_gauss_blur_2_update_0_stage_177 <= dark_gauss_blur_2_update_0_stage_176;
      dark_gauss_blur_2_update_0_stage_178 <= dark_gauss_blur_2_update_0_stage_177;
      dark_gauss_blur_2_update_0_stage_179 <= dark_gauss_blur_2_update_0_stage_178;
      dark_gauss_blur_2_update_0_stage_180 <= dark_gauss_blur_2_update_0_stage_179;
      dark_gauss_blur_2_update_0_stage_181 <= dark_gauss_blur_2_update_0_stage_180;
      bright_gauss_ds_1_update_0_stage_33 <= bright_gauss_ds_1_update_0;
      bright_gauss_ds_1_update_0_stage_34 <= bright_gauss_ds_1_update_0_stage_33;
      bright_gauss_ds_1_update_0_stage_35 <= bright_gauss_ds_1_update_0_stage_34;
      bright_gauss_ds_1_update_0_stage_36 <= bright_gauss_ds_1_update_0_stage_35;
      bright_gauss_ds_1_update_0_stage_37 <= bright_gauss_ds_1_update_0_stage_36;
      bright_gauss_ds_1_update_0_stage_38 <= bright_gauss_ds_1_update_0_stage_37;
      bright_gauss_ds_1_update_0_stage_39 <= bright_gauss_ds_1_update_0_stage_38;
      bright_gauss_ds_1_update_0_stage_40 <= bright_gauss_ds_1_update_0_stage_39;
      bright_gauss_ds_1_update_0_stage_41 <= bright_gauss_ds_1_update_0_stage_40;
      bright_gauss_ds_1_update_0_stage_42 <= bright_gauss_ds_1_update_0_stage_41;
      bright_gauss_ds_1_update_0_stage_43 <= bright_gauss_ds_1_update_0_stage_42;
      bright_gauss_ds_1_update_0_stage_44 <= bright_gauss_ds_1_update_0_stage_43;
      bright_gauss_ds_1_update_0_stage_45 <= bright_gauss_ds_1_update_0_stage_44;
      bright_gauss_ds_1_update_0_stage_46 <= bright_gauss_ds_1_update_0_stage_45;
      bright_gauss_ds_1_update_0_stage_47 <= bright_gauss_ds_1_update_0_stage_46;
      bright_gauss_ds_1_update_0_stage_48 <= bright_gauss_ds_1_update_0_stage_47;
      bright_gauss_ds_1_update_0_stage_49 <= bright_gauss_ds_1_update_0_stage_48;
      bright_gauss_ds_1_update_0_stage_50 <= bright_gauss_ds_1_update_0_stage_49;
      bright_gauss_ds_1_update_0_stage_51 <= bright_gauss_ds_1_update_0_stage_50;
      bright_gauss_ds_1_update_0_stage_52 <= bright_gauss_ds_1_update_0_stage_51;
      bright_gauss_ds_1_update_0_stage_53 <= bright_gauss_ds_1_update_0_stage_52;
      bright_gauss_ds_1_update_0_stage_54 <= bright_gauss_ds_1_update_0_stage_53;
      bright_gauss_ds_1_update_0_stage_55 <= bright_gauss_ds_1_update_0_stage_54;
      bright_gauss_ds_1_update_0_stage_56 <= bright_gauss_ds_1_update_0_stage_55;
      bright_gauss_ds_1_update_0_stage_57 <= bright_gauss_ds_1_update_0_stage_56;
      bright_gauss_ds_1_update_0_stage_58 <= bright_gauss_ds_1_update_0_stage_57;
      bright_gauss_ds_1_update_0_stage_59 <= bright_gauss_ds_1_update_0_stage_58;
      bright_gauss_ds_1_update_0_stage_60 <= bright_gauss_ds_1_update_0_stage_59;
      bright_gauss_ds_1_update_0_stage_61 <= bright_gauss_ds_1_update_0_stage_60;
      bright_gauss_ds_1_update_0_stage_62 <= bright_gauss_ds_1_update_0_stage_61;
      bright_gauss_ds_1_update_0_stage_63 <= bright_gauss_ds_1_update_0_stage_62;
      bright_gauss_ds_1_update_0_stage_64 <= bright_gauss_ds_1_update_0_stage_63;
      bright_gauss_ds_1_update_0_stage_65 <= bright_gauss_ds_1_update_0_stage_64;
      bright_gauss_ds_1_update_0_stage_66 <= bright_gauss_ds_1_update_0_stage_65;
      bright_gauss_ds_1_update_0_stage_67 <= bright_gauss_ds_1_update_0_stage_66;
      bright_gauss_ds_1_update_0_stage_68 <= bright_gauss_ds_1_update_0_stage_67;
      bright_gauss_ds_1_update_0_stage_69 <= bright_gauss_ds_1_update_0_stage_68;
      bright_gauss_ds_1_update_0_stage_70 <= bright_gauss_ds_1_update_0_stage_69;
      bright_gauss_ds_1_update_0_stage_71 <= bright_gauss_ds_1_update_0_stage_70;
      bright_gauss_ds_1_update_0_stage_72 <= bright_gauss_ds_1_update_0_stage_71;
      bright_gauss_ds_1_update_0_stage_73 <= bright_gauss_ds_1_update_0_stage_72;
      bright_gauss_ds_1_update_0_stage_74 <= bright_gauss_ds_1_update_0_stage_73;
      bright_gauss_ds_1_update_0_stage_75 <= bright_gauss_ds_1_update_0_stage_74;
      bright_gauss_ds_1_update_0_stage_76 <= bright_gauss_ds_1_update_0_stage_75;
      bright_gauss_ds_1_update_0_stage_77 <= bright_gauss_ds_1_update_0_stage_76;
      bright_gauss_ds_1_update_0_stage_78 <= bright_gauss_ds_1_update_0_stage_77;
      bright_gauss_ds_1_update_0_stage_79 <= bright_gauss_ds_1_update_0_stage_78;
      bright_gauss_ds_1_update_0_stage_80 <= bright_gauss_ds_1_update_0_stage_79;
      bright_gauss_ds_1_update_0_stage_81 <= bright_gauss_ds_1_update_0_stage_80;
      bright_gauss_ds_1_update_0_stage_82 <= bright_gauss_ds_1_update_0_stage_81;
      bright_gauss_ds_1_update_0_stage_83 <= bright_gauss_ds_1_update_0_stage_82;
      bright_gauss_ds_1_update_0_stage_84 <= bright_gauss_ds_1_update_0_stage_83;
      bright_gauss_ds_1_update_0_stage_85 <= bright_gauss_ds_1_update_0_stage_84;
      bright_gauss_ds_1_update_0_stage_86 <= bright_gauss_ds_1_update_0_stage_85;
      bright_gauss_ds_1_update_0_stage_87 <= bright_gauss_ds_1_update_0_stage_86;
      bright_gauss_ds_1_update_0_stage_88 <= bright_gauss_ds_1_update_0_stage_87;
      bright_gauss_ds_1_update_0_stage_89 <= bright_gauss_ds_1_update_0_stage_88;
      bright_gauss_ds_1_update_0_stage_90 <= bright_gauss_ds_1_update_0_stage_89;
      bright_gauss_ds_1_update_0_stage_91 <= bright_gauss_ds_1_update_0_stage_90;
      bright_gauss_ds_1_update_0_stage_92 <= bright_gauss_ds_1_update_0_stage_91;
      bright_gauss_ds_1_update_0_stage_93 <= bright_gauss_ds_1_update_0_stage_92;
      bright_gauss_ds_1_update_0_stage_94 <= bright_gauss_ds_1_update_0_stage_93;
      bright_gauss_ds_1_update_0_stage_95 <= bright_gauss_ds_1_update_0_stage_94;
      bright_gauss_ds_1_update_0_stage_96 <= bright_gauss_ds_1_update_0_stage_95;
      bright_gauss_ds_1_update_0_stage_97 <= bright_gauss_ds_1_update_0_stage_96;
      bright_gauss_ds_1_update_0_stage_98 <= bright_gauss_ds_1_update_0_stage_97;
      bright_gauss_ds_1_update_0_stage_99 <= bright_gauss_ds_1_update_0_stage_98;
      bright_gauss_ds_1_update_0_stage_100 <= bright_gauss_ds_1_update_0_stage_99;
      bright_gauss_ds_1_update_0_stage_101 <= bright_gauss_ds_1_update_0_stage_100;
      bright_gauss_ds_1_update_0_stage_102 <= bright_gauss_ds_1_update_0_stage_101;
      bright_gauss_ds_1_update_0_stage_103 <= bright_gauss_ds_1_update_0_stage_102;
      bright_gauss_ds_1_update_0_stage_104 <= bright_gauss_ds_1_update_0_stage_103;
      bright_gauss_ds_1_update_0_stage_105 <= bright_gauss_ds_1_update_0_stage_104;
      bright_gauss_ds_1_update_0_stage_106 <= bright_gauss_ds_1_update_0_stage_105;
      bright_gauss_ds_1_update_0_stage_107 <= bright_gauss_ds_1_update_0_stage_106;
      bright_gauss_ds_1_update_0_stage_108 <= bright_gauss_ds_1_update_0_stage_107;
      bright_gauss_ds_1_update_0_stage_109 <= bright_gauss_ds_1_update_0_stage_108;
      bright_gauss_ds_1_update_0_stage_110 <= bright_gauss_ds_1_update_0_stage_109;
      bright_gauss_ds_1_update_0_stage_111 <= bright_gauss_ds_1_update_0_stage_110;
      bright_gauss_ds_1_update_0_stage_112 <= bright_gauss_ds_1_update_0_stage_111;
      bright_gauss_ds_1_update_0_stage_113 <= bright_gauss_ds_1_update_0_stage_112;
      bright_gauss_ds_1_update_0_stage_114 <= bright_gauss_ds_1_update_0_stage_113;
      bright_gauss_ds_1_update_0_stage_115 <= bright_gauss_ds_1_update_0_stage_114;
      bright_gauss_ds_1_update_0_stage_116 <= bright_gauss_ds_1_update_0_stage_115;
      bright_gauss_ds_1_update_0_stage_117 <= bright_gauss_ds_1_update_0_stage_116;
      bright_gauss_ds_1_update_0_stage_118 <= bright_gauss_ds_1_update_0_stage_117;
      bright_gauss_ds_1_update_0_stage_119 <= bright_gauss_ds_1_update_0_stage_118;
      bright_gauss_ds_1_update_0_stage_120 <= bright_gauss_ds_1_update_0_stage_119;
      bright_gauss_ds_1_update_0_stage_121 <= bright_gauss_ds_1_update_0_stage_120;
      bright_gauss_ds_1_update_0_stage_122 <= bright_gauss_ds_1_update_0_stage_121;
      bright_gauss_ds_1_update_0_stage_123 <= bright_gauss_ds_1_update_0_stage_122;
      bright_gauss_ds_1_update_0_stage_124 <= bright_gauss_ds_1_update_0_stage_123;
      bright_gauss_ds_1_update_0_stage_125 <= bright_gauss_ds_1_update_0_stage_124;
      bright_gauss_ds_1_update_0_stage_126 <= bright_gauss_ds_1_update_0_stage_125;
      bright_gauss_ds_1_update_0_stage_127 <= bright_gauss_ds_1_update_0_stage_126;
      bright_gauss_ds_1_update_0_stage_128 <= bright_gauss_ds_1_update_0_stage_127;
      bright_gauss_ds_1_update_0_stage_129 <= bright_gauss_ds_1_update_0_stage_128;
      bright_gauss_ds_1_update_0_stage_130 <= bright_gauss_ds_1_update_0_stage_129;
      bright_gauss_ds_1_update_0_stage_131 <= bright_gauss_ds_1_update_0_stage_130;
      bright_gauss_ds_1_update_0_stage_132 <= bright_gauss_ds_1_update_0_stage_131;
      bright_gauss_ds_1_update_0_stage_133 <= bright_gauss_ds_1_update_0_stage_132;
      bright_gauss_ds_1_update_0_stage_134 <= bright_gauss_ds_1_update_0_stage_133;
      bright_gauss_ds_1_update_0_stage_135 <= bright_gauss_ds_1_update_0_stage_134;
      bright_gauss_ds_1_update_0_stage_136 <= bright_gauss_ds_1_update_0_stage_135;
      bright_gauss_ds_1_update_0_stage_137 <= bright_gauss_ds_1_update_0_stage_136;
      bright_gauss_ds_1_update_0_stage_138 <= bright_gauss_ds_1_update_0_stage_137;
      bright_gauss_ds_1_update_0_stage_139 <= bright_gauss_ds_1_update_0_stage_138;
      bright_gauss_ds_1_update_0_stage_140 <= bright_gauss_ds_1_update_0_stage_139;
      bright_gauss_ds_1_update_0_stage_141 <= bright_gauss_ds_1_update_0_stage_140;
      bright_gauss_ds_1_update_0_stage_142 <= bright_gauss_ds_1_update_0_stage_141;
      bright_gauss_ds_1_update_0_stage_143 <= bright_gauss_ds_1_update_0_stage_142;
      bright_gauss_ds_1_update_0_stage_144 <= bright_gauss_ds_1_update_0_stage_143;
      bright_gauss_ds_1_update_0_stage_145 <= bright_gauss_ds_1_update_0_stage_144;
      bright_gauss_ds_1_update_0_stage_146 <= bright_gauss_ds_1_update_0_stage_145;
      bright_gauss_ds_1_update_0_stage_147 <= bright_gauss_ds_1_update_0_stage_146;
      bright_gauss_ds_1_update_0_stage_148 <= bright_gauss_ds_1_update_0_stage_147;
      bright_gauss_ds_1_update_0_stage_149 <= bright_gauss_ds_1_update_0_stage_148;
      bright_gauss_ds_1_update_0_stage_150 <= bright_gauss_ds_1_update_0_stage_149;
      bright_gauss_ds_1_update_0_stage_151 <= bright_gauss_ds_1_update_0_stage_150;
      bright_gauss_ds_1_update_0_stage_152 <= bright_gauss_ds_1_update_0_stage_151;
      bright_gauss_ds_1_update_0_stage_153 <= bright_gauss_ds_1_update_0_stage_152;
      bright_gauss_ds_1_update_0_stage_154 <= bright_gauss_ds_1_update_0_stage_153;
      bright_gauss_ds_1_update_0_stage_155 <= bright_gauss_ds_1_update_0_stage_154;
      bright_gauss_ds_1_update_0_stage_156 <= bright_gauss_ds_1_update_0_stage_155;
      bright_gauss_ds_1_update_0_stage_157 <= bright_gauss_ds_1_update_0_stage_156;
      bright_gauss_ds_1_update_0_stage_158 <= bright_gauss_ds_1_update_0_stage_157;
      bright_gauss_ds_1_update_0_stage_159 <= bright_gauss_ds_1_update_0_stage_158;
      bright_gauss_ds_1_update_0_stage_160 <= bright_gauss_ds_1_update_0_stage_159;
      bright_gauss_ds_1_update_0_stage_161 <= bright_gauss_ds_1_update_0_stage_160;
      bright_gauss_ds_1_update_0_stage_162 <= bright_gauss_ds_1_update_0_stage_161;
      bright_gauss_ds_1_update_0_stage_163 <= bright_gauss_ds_1_update_0_stage_162;
      bright_gauss_ds_1_update_0_stage_164 <= bright_gauss_ds_1_update_0_stage_163;
      bright_gauss_ds_1_update_0_stage_165 <= bright_gauss_ds_1_update_0_stage_164;
      bright_gauss_ds_1_update_0_stage_166 <= bright_gauss_ds_1_update_0_stage_165;
      bright_gauss_ds_1_update_0_stage_167 <= bright_gauss_ds_1_update_0_stage_166;
      bright_gauss_ds_1_update_0_stage_168 <= bright_gauss_ds_1_update_0_stage_167;
      bright_gauss_ds_1_update_0_stage_169 <= bright_gauss_ds_1_update_0_stage_168;
      bright_gauss_ds_1_update_0_stage_170 <= bright_gauss_ds_1_update_0_stage_169;
      bright_gauss_ds_1_update_0_stage_171 <= bright_gauss_ds_1_update_0_stage_170;
      bright_gauss_ds_1_update_0_stage_172 <= bright_gauss_ds_1_update_0_stage_171;
      bright_gauss_ds_1_update_0_stage_173 <= bright_gauss_ds_1_update_0_stage_172;
      bright_gauss_ds_1_update_0_stage_174 <= bright_gauss_ds_1_update_0_stage_173;
      bright_gauss_ds_1_update_0_stage_175 <= bright_gauss_ds_1_update_0_stage_174;
      bright_gauss_ds_1_update_0_stage_176 <= bright_gauss_ds_1_update_0_stage_175;
      bright_gauss_ds_1_update_0_stage_177 <= bright_gauss_ds_1_update_0_stage_176;
      bright_gauss_ds_1_update_0_stage_178 <= bright_gauss_ds_1_update_0_stage_177;
      bright_gauss_ds_1_update_0_stage_179 <= bright_gauss_ds_1_update_0_stage_178;
      bright_gauss_ds_1_update_0_stage_180 <= bright_gauss_ds_1_update_0_stage_179;
      bright_gauss_ds_1_update_0_stage_181 <= bright_gauss_ds_1_update_0_stage_180;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_34 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_35 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_34;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_36 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_35;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_37 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_36;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_38 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_37;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_39 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_38;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_40 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_39;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_41 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_40;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_42 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_41;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_43 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_42;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_44 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_43;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_45 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_44;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_46 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_45;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_47 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_46;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_48 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_47;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_49 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_48;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_50 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_49;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_51 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_50;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_52 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_51;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_53 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_52;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_54 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_53;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_55 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_54;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_56 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_55;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_57 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_56;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_58 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_57;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_59 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_58;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_60 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_59;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_61 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_60;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_62 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_61;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_63 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_62;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_64 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_63;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_65 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_64;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_66 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_65;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_67 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_66;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_68 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_67;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_69 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_68;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_70 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_69;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_71 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_70;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_72 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_71;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_73 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_72;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_74 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_73;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_75 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_74;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_76 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_75;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_77 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_76;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_78 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_77;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_79 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_78;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_80 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_79;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_81 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_80;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_82 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_81;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_83 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_82;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_84 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_83;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_85 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_84;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_86 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_85;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_87 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_86;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_88 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_87;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_89 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_88;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_90 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_89;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_91 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_90;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_92 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_91;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_93 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_92;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_94 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_93;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_95 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_94;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_96 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_95;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_97 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_96;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_98 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_97;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_99 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_98;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_100 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_99;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_101 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_100;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_102 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_101;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_103 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_102;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_104 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_103;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_105 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_104;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_106 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_105;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_107 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_106;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_108 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_107;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_109 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_108;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_110 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_109;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_111 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_110;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_112 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_111;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_113 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_112;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_114 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_113;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_115 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_114;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_116 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_115;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_117 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_116;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_118 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_117;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_119 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_118;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_120 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_119;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_121 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_120;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_122 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_121;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_123 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_122;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_124 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_123;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_125 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_124;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_126 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_125;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_127 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_126;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_128 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_127;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_129 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_128;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_130 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_129;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_131 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_130;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_132 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_131;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_133 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_132;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_134 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_133;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_135 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_134;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_136 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_135;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_137 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_136;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_138 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_137;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_139 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_138;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_140 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_139;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_141 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_140;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_142 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_141;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_143 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_142;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_144 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_143;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_145 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_144;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_146 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_145;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_147 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_146;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_148 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_147;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_149 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_148;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_150 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_149;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_151 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_150;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_152 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_151;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_153 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_152;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_154 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_153;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_155 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_154;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_156 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_155;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_157 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_156;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_158 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_157;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_159 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_158;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_160 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_159;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_161 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_160;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_162 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_161;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_163 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_162;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_164 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_163;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_165 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_164;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_166 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_165;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_167 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_166;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_168 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_167;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_169 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_168;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_170 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_169;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_171 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_170;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_172 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_171;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_173 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_172;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_174 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_173;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_175 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_174;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_176 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_175;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_177 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_176;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_178 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_177;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_179 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_178;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_180 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_179;
      bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_181 <= bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21_stage_180;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_69 <= weight_sums_dark_weights_normed_update_0_read_read_46;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_70 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_69;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_71 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_70;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_72 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_71;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_73 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_72;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_74 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_73;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_75 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_74;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_76 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_75;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_77 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_76;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_78 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_77;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_79 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_78;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_80 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_79;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_81 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_80;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_82 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_81;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_83 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_82;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_84 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_83;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_85 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_84;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_86 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_85;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_87 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_86;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_88 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_87;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_89 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_88;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_90 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_89;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_91 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_90;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_92 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_91;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_93 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_92;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_94 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_93;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_95 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_94;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_96 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_95;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_97 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_96;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_98 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_97;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_99 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_98;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_100 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_99;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_101 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_100;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_102 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_101;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_103 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_102;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_104 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_103;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_105 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_104;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_106 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_105;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_107 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_106;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_108 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_107;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_109 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_108;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_110 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_109;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_111 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_110;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_112 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_111;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_113 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_112;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_114 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_113;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_115 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_114;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_116 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_115;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_117 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_116;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_118 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_117;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_119 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_118;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_120 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_119;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_121 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_120;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_122 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_121;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_123 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_122;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_124 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_123;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_125 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_124;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_126 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_125;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_127 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_126;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_128 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_127;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_129 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_128;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_130 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_129;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_131 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_130;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_132 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_131;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_133 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_132;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_134 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_133;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_135 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_134;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_136 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_135;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_137 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_136;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_138 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_137;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_139 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_138;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_140 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_139;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_141 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_140;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_142 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_141;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_143 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_142;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_144 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_143;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_145 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_144;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_146 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_145;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_147 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_146;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_148 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_147;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_149 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_148;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_150 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_149;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_151 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_150;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_152 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_151;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_153 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_152;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_154 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_153;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_155 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_154;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_156 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_155;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_157 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_156;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_158 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_157;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_159 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_158;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_160 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_159;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_161 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_160;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_162 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_161;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_163 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_162;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_164 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_163;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_165 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_164;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_166 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_165;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_167 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_166;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_168 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_167;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_169 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_168;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_170 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_169;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_171 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_170;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_172 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_171;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_173 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_172;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_174 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_173;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_175 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_174;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_176 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_175;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_177 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_176;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_178 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_177;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_179 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_178;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_180 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_179;
      weight_sums_dark_weights_normed_update_0_read_read_46_stage_181 <= weight_sums_dark_weights_normed_update_0_read_read_46_stage_180;
      dark_weights_normed_update_0_stage_70 <= dark_weights_normed_update_0;
      dark_weights_normed_update_0_stage_71 <= dark_weights_normed_update_0_stage_70;
      dark_weights_normed_update_0_stage_72 <= dark_weights_normed_update_0_stage_71;
      dark_weights_normed_update_0_stage_73 <= dark_weights_normed_update_0_stage_72;
      dark_weights_normed_update_0_stage_74 <= dark_weights_normed_update_0_stage_73;
      dark_weights_normed_update_0_stage_75 <= dark_weights_normed_update_0_stage_74;
      dark_weights_normed_update_0_stage_76 <= dark_weights_normed_update_0_stage_75;
      dark_weights_normed_update_0_stage_77 <= dark_weights_normed_update_0_stage_76;
      dark_weights_normed_update_0_stage_78 <= dark_weights_normed_update_0_stage_77;
      dark_weights_normed_update_0_stage_79 <= dark_weights_normed_update_0_stage_78;
      dark_weights_normed_update_0_stage_80 <= dark_weights_normed_update_0_stage_79;
      dark_weights_normed_update_0_stage_81 <= dark_weights_normed_update_0_stage_80;
      dark_weights_normed_update_0_stage_82 <= dark_weights_normed_update_0_stage_81;
      dark_weights_normed_update_0_stage_83 <= dark_weights_normed_update_0_stage_82;
      dark_weights_normed_update_0_stage_84 <= dark_weights_normed_update_0_stage_83;
      dark_weights_normed_update_0_stage_85 <= dark_weights_normed_update_0_stage_84;
      dark_weights_normed_update_0_stage_86 <= dark_weights_normed_update_0_stage_85;
      dark_weights_normed_update_0_stage_87 <= dark_weights_normed_update_0_stage_86;
      dark_weights_normed_update_0_stage_88 <= dark_weights_normed_update_0_stage_87;
      dark_weights_normed_update_0_stage_89 <= dark_weights_normed_update_0_stage_88;
      dark_weights_normed_update_0_stage_90 <= dark_weights_normed_update_0_stage_89;
      dark_weights_normed_update_0_stage_91 <= dark_weights_normed_update_0_stage_90;
      dark_weights_normed_update_0_stage_92 <= dark_weights_normed_update_0_stage_91;
      dark_weights_normed_update_0_stage_93 <= dark_weights_normed_update_0_stage_92;
      dark_weights_normed_update_0_stage_94 <= dark_weights_normed_update_0_stage_93;
      dark_weights_normed_update_0_stage_95 <= dark_weights_normed_update_0_stage_94;
      dark_weights_normed_update_0_stage_96 <= dark_weights_normed_update_0_stage_95;
      dark_weights_normed_update_0_stage_97 <= dark_weights_normed_update_0_stage_96;
      dark_weights_normed_update_0_stage_98 <= dark_weights_normed_update_0_stage_97;
      dark_weights_normed_update_0_stage_99 <= dark_weights_normed_update_0_stage_98;
      dark_weights_normed_update_0_stage_100 <= dark_weights_normed_update_0_stage_99;
      dark_weights_normed_update_0_stage_101 <= dark_weights_normed_update_0_stage_100;
      dark_weights_normed_update_0_stage_102 <= dark_weights_normed_update_0_stage_101;
      dark_weights_normed_update_0_stage_103 <= dark_weights_normed_update_0_stage_102;
      dark_weights_normed_update_0_stage_104 <= dark_weights_normed_update_0_stage_103;
      dark_weights_normed_update_0_stage_105 <= dark_weights_normed_update_0_stage_104;
      dark_weights_normed_update_0_stage_106 <= dark_weights_normed_update_0_stage_105;
      dark_weights_normed_update_0_stage_107 <= dark_weights_normed_update_0_stage_106;
      dark_weights_normed_update_0_stage_108 <= dark_weights_normed_update_0_stage_107;
      dark_weights_normed_update_0_stage_109 <= dark_weights_normed_update_0_stage_108;
      dark_weights_normed_update_0_stage_110 <= dark_weights_normed_update_0_stage_109;
      dark_weights_normed_update_0_stage_111 <= dark_weights_normed_update_0_stage_110;
      dark_weights_normed_update_0_stage_112 <= dark_weights_normed_update_0_stage_111;
      dark_weights_normed_update_0_stage_113 <= dark_weights_normed_update_0_stage_112;
      dark_weights_normed_update_0_stage_114 <= dark_weights_normed_update_0_stage_113;
      dark_weights_normed_update_0_stage_115 <= dark_weights_normed_update_0_stage_114;
      dark_weights_normed_update_0_stage_116 <= dark_weights_normed_update_0_stage_115;
      dark_weights_normed_update_0_stage_117 <= dark_weights_normed_update_0_stage_116;
      dark_weights_normed_update_0_stage_118 <= dark_weights_normed_update_0_stage_117;
      dark_weights_normed_update_0_stage_119 <= dark_weights_normed_update_0_stage_118;
      dark_weights_normed_update_0_stage_120 <= dark_weights_normed_update_0_stage_119;
      dark_weights_normed_update_0_stage_121 <= dark_weights_normed_update_0_stage_120;
      dark_weights_normed_update_0_stage_122 <= dark_weights_normed_update_0_stage_121;
      dark_weights_normed_update_0_stage_123 <= dark_weights_normed_update_0_stage_122;
      dark_weights_normed_update_0_stage_124 <= dark_weights_normed_update_0_stage_123;
      dark_weights_normed_update_0_stage_125 <= dark_weights_normed_update_0_stage_124;
      dark_weights_normed_update_0_stage_126 <= dark_weights_normed_update_0_stage_125;
      dark_weights_normed_update_0_stage_127 <= dark_weights_normed_update_0_stage_126;
      dark_weights_normed_update_0_stage_128 <= dark_weights_normed_update_0_stage_127;
      dark_weights_normed_update_0_stage_129 <= dark_weights_normed_update_0_stage_128;
      dark_weights_normed_update_0_stage_130 <= dark_weights_normed_update_0_stage_129;
      dark_weights_normed_update_0_stage_131 <= dark_weights_normed_update_0_stage_130;
      dark_weights_normed_update_0_stage_132 <= dark_weights_normed_update_0_stage_131;
      dark_weights_normed_update_0_stage_133 <= dark_weights_normed_update_0_stage_132;
      dark_weights_normed_update_0_stage_134 <= dark_weights_normed_update_0_stage_133;
      dark_weights_normed_update_0_stage_135 <= dark_weights_normed_update_0_stage_134;
      dark_weights_normed_update_0_stage_136 <= dark_weights_normed_update_0_stage_135;
      dark_weights_normed_update_0_stage_137 <= dark_weights_normed_update_0_stage_136;
      dark_weights_normed_update_0_stage_138 <= dark_weights_normed_update_0_stage_137;
      dark_weights_normed_update_0_stage_139 <= dark_weights_normed_update_0_stage_138;
      dark_weights_normed_update_0_stage_140 <= dark_weights_normed_update_0_stage_139;
      dark_weights_normed_update_0_stage_141 <= dark_weights_normed_update_0_stage_140;
      dark_weights_normed_update_0_stage_142 <= dark_weights_normed_update_0_stage_141;
      dark_weights_normed_update_0_stage_143 <= dark_weights_normed_update_0_stage_142;
      dark_weights_normed_update_0_stage_144 <= dark_weights_normed_update_0_stage_143;
      dark_weights_normed_update_0_stage_145 <= dark_weights_normed_update_0_stage_144;
      dark_weights_normed_update_0_stage_146 <= dark_weights_normed_update_0_stage_145;
      dark_weights_normed_update_0_stage_147 <= dark_weights_normed_update_0_stage_146;
      dark_weights_normed_update_0_stage_148 <= dark_weights_normed_update_0_stage_147;
      dark_weights_normed_update_0_stage_149 <= dark_weights_normed_update_0_stage_148;
      dark_weights_normed_update_0_stage_150 <= dark_weights_normed_update_0_stage_149;
      dark_weights_normed_update_0_stage_151 <= dark_weights_normed_update_0_stage_150;
      dark_weights_normed_update_0_stage_152 <= dark_weights_normed_update_0_stage_151;
      dark_weights_normed_update_0_stage_153 <= dark_weights_normed_update_0_stage_152;
      dark_weights_normed_update_0_stage_154 <= dark_weights_normed_update_0_stage_153;
      dark_weights_normed_update_0_stage_155 <= dark_weights_normed_update_0_stage_154;
      dark_weights_normed_update_0_stage_156 <= dark_weights_normed_update_0_stage_155;
      dark_weights_normed_update_0_stage_157 <= dark_weights_normed_update_0_stage_156;
      dark_weights_normed_update_0_stage_158 <= dark_weights_normed_update_0_stage_157;
      dark_weights_normed_update_0_stage_159 <= dark_weights_normed_update_0_stage_158;
      dark_weights_normed_update_0_stage_160 <= dark_weights_normed_update_0_stage_159;
      dark_weights_normed_update_0_stage_161 <= dark_weights_normed_update_0_stage_160;
      dark_weights_normed_update_0_stage_162 <= dark_weights_normed_update_0_stage_161;
      dark_weights_normed_update_0_stage_163 <= dark_weights_normed_update_0_stage_162;
      dark_weights_normed_update_0_stage_164 <= dark_weights_normed_update_0_stage_163;
      dark_weights_normed_update_0_stage_165 <= dark_weights_normed_update_0_stage_164;
      dark_weights_normed_update_0_stage_166 <= dark_weights_normed_update_0_stage_165;
      dark_weights_normed_update_0_stage_167 <= dark_weights_normed_update_0_stage_166;
      dark_weights_normed_update_0_stage_168 <= dark_weights_normed_update_0_stage_167;
      dark_weights_normed_update_0_stage_169 <= dark_weights_normed_update_0_stage_168;
      dark_weights_normed_update_0_stage_170 <= dark_weights_normed_update_0_stage_169;
      dark_weights_normed_update_0_stage_171 <= dark_weights_normed_update_0_stage_170;
      dark_weights_normed_update_0_stage_172 <= dark_weights_normed_update_0_stage_171;
      dark_weights_normed_update_0_stage_173 <= dark_weights_normed_update_0_stage_172;
      dark_weights_normed_update_0_stage_174 <= dark_weights_normed_update_0_stage_173;
      dark_weights_normed_update_0_stage_175 <= dark_weights_normed_update_0_stage_174;
      dark_weights_normed_update_0_stage_176 <= dark_weights_normed_update_0_stage_175;
      dark_weights_normed_update_0_stage_177 <= dark_weights_normed_update_0_stage_176;
      dark_weights_normed_update_0_stage_178 <= dark_weights_normed_update_0_stage_177;
      dark_weights_normed_update_0_stage_179 <= dark_weights_normed_update_0_stage_178;
      dark_weights_normed_update_0_stage_180 <= dark_weights_normed_update_0_stage_179;
      dark_weights_normed_update_0_stage_181 <= dark_weights_normed_update_0_stage_180;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_39 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_40 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_39;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_41 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_40;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_42 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_41;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_43 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_42;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_44 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_43;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_45 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_44;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_46 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_45;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_47 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_46;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_48 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_47;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_49 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_48;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_50 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_49;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_51 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_50;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_52 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_51;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_53 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_52;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_54 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_53;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_55 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_54;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_56 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_55;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_57 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_56;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_58 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_57;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_59 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_58;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_60 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_59;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_61 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_60;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_62 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_61;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_63 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_62;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_64 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_63;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_65 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_64;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_66 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_65;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_67 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_66;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_68 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_67;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_69 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_68;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_70 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_69;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_71 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_70;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_72 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_71;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_73 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_72;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_74 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_73;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_75 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_74;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_76 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_75;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_77 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_76;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_78 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_77;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_79 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_78;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_80 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_79;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_81 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_80;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_82 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_81;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_83 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_82;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_84 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_83;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_85 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_84;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_86 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_85;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_87 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_86;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_88 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_87;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_89 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_88;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_90 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_89;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_91 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_90;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_92 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_91;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_93 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_92;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_94 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_93;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_95 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_94;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_96 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_95;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_97 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_96;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_98 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_97;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_99 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_98;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_100 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_99;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_101 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_100;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_102 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_101;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_103 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_102;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_104 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_103;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_105 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_104;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_106 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_105;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_107 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_106;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_108 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_107;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_109 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_108;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_110 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_109;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_111 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_110;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_112 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_111;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_113 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_112;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_114 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_113;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_115 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_114;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_116 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_115;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_117 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_116;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_118 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_117;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_119 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_118;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_120 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_119;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_121 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_120;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_122 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_121;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_123 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_122;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_124 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_123;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_125 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_124;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_126 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_125;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_127 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_126;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_128 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_127;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_129 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_128;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_130 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_129;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_131 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_130;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_132 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_131;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_133 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_132;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_134 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_133;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_135 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_134;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_136 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_135;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_137 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_136;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_138 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_137;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_139 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_138;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_140 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_139;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_141 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_140;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_142 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_141;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_143 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_142;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_144 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_143;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_145 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_144;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_146 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_145;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_147 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_146;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_148 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_147;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_149 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_148;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_150 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_149;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_151 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_150;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_152 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_151;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_153 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_152;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_154 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_153;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_155 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_154;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_156 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_155;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_157 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_156;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_158 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_157;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_159 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_158;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_160 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_159;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_161 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_160;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_162 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_161;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_163 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_162;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_164 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_163;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_165 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_164;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_166 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_165;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_167 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_166;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_168 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_167;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_169 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_168;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_170 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_169;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_171 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_170;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_172 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_171;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_173 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_172;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_174 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_173;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_175 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_174;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_176 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_175;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_177 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_176;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_178 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_177;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_179 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_178;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_180 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_179;
      bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_181 <= bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25_stage_180;
      bright_gauss_blur_2_update_0_stage_40 <= bright_gauss_blur_2_update_0;
      bright_gauss_blur_2_update_0_stage_41 <= bright_gauss_blur_2_update_0_stage_40;
      bright_gauss_blur_2_update_0_stage_42 <= bright_gauss_blur_2_update_0_stage_41;
      bright_gauss_blur_2_update_0_stage_43 <= bright_gauss_blur_2_update_0_stage_42;
      bright_gauss_blur_2_update_0_stage_44 <= bright_gauss_blur_2_update_0_stage_43;
      bright_gauss_blur_2_update_0_stage_45 <= bright_gauss_blur_2_update_0_stage_44;
      bright_gauss_blur_2_update_0_stage_46 <= bright_gauss_blur_2_update_0_stage_45;
      bright_gauss_blur_2_update_0_stage_47 <= bright_gauss_blur_2_update_0_stage_46;
      bright_gauss_blur_2_update_0_stage_48 <= bright_gauss_blur_2_update_0_stage_47;
      bright_gauss_blur_2_update_0_stage_49 <= bright_gauss_blur_2_update_0_stage_48;
      bright_gauss_blur_2_update_0_stage_50 <= bright_gauss_blur_2_update_0_stage_49;
      bright_gauss_blur_2_update_0_stage_51 <= bright_gauss_blur_2_update_0_stage_50;
      bright_gauss_blur_2_update_0_stage_52 <= bright_gauss_blur_2_update_0_stage_51;
      bright_gauss_blur_2_update_0_stage_53 <= bright_gauss_blur_2_update_0_stage_52;
      bright_gauss_blur_2_update_0_stage_54 <= bright_gauss_blur_2_update_0_stage_53;
      bright_gauss_blur_2_update_0_stage_55 <= bright_gauss_blur_2_update_0_stage_54;
      bright_gauss_blur_2_update_0_stage_56 <= bright_gauss_blur_2_update_0_stage_55;
      bright_gauss_blur_2_update_0_stage_57 <= bright_gauss_blur_2_update_0_stage_56;
      bright_gauss_blur_2_update_0_stage_58 <= bright_gauss_blur_2_update_0_stage_57;
      bright_gauss_blur_2_update_0_stage_59 <= bright_gauss_blur_2_update_0_stage_58;
      bright_gauss_blur_2_update_0_stage_60 <= bright_gauss_blur_2_update_0_stage_59;
      bright_gauss_blur_2_update_0_stage_61 <= bright_gauss_blur_2_update_0_stage_60;
      bright_gauss_blur_2_update_0_stage_62 <= bright_gauss_blur_2_update_0_stage_61;
      bright_gauss_blur_2_update_0_stage_63 <= bright_gauss_blur_2_update_0_stage_62;
      bright_gauss_blur_2_update_0_stage_64 <= bright_gauss_blur_2_update_0_stage_63;
      bright_gauss_blur_2_update_0_stage_65 <= bright_gauss_blur_2_update_0_stage_64;
      bright_gauss_blur_2_update_0_stage_66 <= bright_gauss_blur_2_update_0_stage_65;
      bright_gauss_blur_2_update_0_stage_67 <= bright_gauss_blur_2_update_0_stage_66;
      bright_gauss_blur_2_update_0_stage_68 <= bright_gauss_blur_2_update_0_stage_67;
      bright_gauss_blur_2_update_0_stage_69 <= bright_gauss_blur_2_update_0_stage_68;
      bright_gauss_blur_2_update_0_stage_70 <= bright_gauss_blur_2_update_0_stage_69;
      bright_gauss_blur_2_update_0_stage_71 <= bright_gauss_blur_2_update_0_stage_70;
      bright_gauss_blur_2_update_0_stage_72 <= bright_gauss_blur_2_update_0_stage_71;
      bright_gauss_blur_2_update_0_stage_73 <= bright_gauss_blur_2_update_0_stage_72;
      bright_gauss_blur_2_update_0_stage_74 <= bright_gauss_blur_2_update_0_stage_73;
      bright_gauss_blur_2_update_0_stage_75 <= bright_gauss_blur_2_update_0_stage_74;
      bright_gauss_blur_2_update_0_stage_76 <= bright_gauss_blur_2_update_0_stage_75;
      bright_gauss_blur_2_update_0_stage_77 <= bright_gauss_blur_2_update_0_stage_76;
      bright_gauss_blur_2_update_0_stage_78 <= bright_gauss_blur_2_update_0_stage_77;
      bright_gauss_blur_2_update_0_stage_79 <= bright_gauss_blur_2_update_0_stage_78;
      bright_gauss_blur_2_update_0_stage_80 <= bright_gauss_blur_2_update_0_stage_79;
      bright_gauss_blur_2_update_0_stage_81 <= bright_gauss_blur_2_update_0_stage_80;
      bright_gauss_blur_2_update_0_stage_82 <= bright_gauss_blur_2_update_0_stage_81;
      bright_gauss_blur_2_update_0_stage_83 <= bright_gauss_blur_2_update_0_stage_82;
      bright_gauss_blur_2_update_0_stage_84 <= bright_gauss_blur_2_update_0_stage_83;
      bright_gauss_blur_2_update_0_stage_85 <= bright_gauss_blur_2_update_0_stage_84;
      bright_gauss_blur_2_update_0_stage_86 <= bright_gauss_blur_2_update_0_stage_85;
      bright_gauss_blur_2_update_0_stage_87 <= bright_gauss_blur_2_update_0_stage_86;
      bright_gauss_blur_2_update_0_stage_88 <= bright_gauss_blur_2_update_0_stage_87;
      bright_gauss_blur_2_update_0_stage_89 <= bright_gauss_blur_2_update_0_stage_88;
      bright_gauss_blur_2_update_0_stage_90 <= bright_gauss_blur_2_update_0_stage_89;
      bright_gauss_blur_2_update_0_stage_91 <= bright_gauss_blur_2_update_0_stage_90;
      bright_gauss_blur_2_update_0_stage_92 <= bright_gauss_blur_2_update_0_stage_91;
      bright_gauss_blur_2_update_0_stage_93 <= bright_gauss_blur_2_update_0_stage_92;
      bright_gauss_blur_2_update_0_stage_94 <= bright_gauss_blur_2_update_0_stage_93;
      bright_gauss_blur_2_update_0_stage_95 <= bright_gauss_blur_2_update_0_stage_94;
      bright_gauss_blur_2_update_0_stage_96 <= bright_gauss_blur_2_update_0_stage_95;
      bright_gauss_blur_2_update_0_stage_97 <= bright_gauss_blur_2_update_0_stage_96;
      bright_gauss_blur_2_update_0_stage_98 <= bright_gauss_blur_2_update_0_stage_97;
      bright_gauss_blur_2_update_0_stage_99 <= bright_gauss_blur_2_update_0_stage_98;
      bright_gauss_blur_2_update_0_stage_100 <= bright_gauss_blur_2_update_0_stage_99;
      bright_gauss_blur_2_update_0_stage_101 <= bright_gauss_blur_2_update_0_stage_100;
      bright_gauss_blur_2_update_0_stage_102 <= bright_gauss_blur_2_update_0_stage_101;
      bright_gauss_blur_2_update_0_stage_103 <= bright_gauss_blur_2_update_0_stage_102;
      bright_gauss_blur_2_update_0_stage_104 <= bright_gauss_blur_2_update_0_stage_103;
      bright_gauss_blur_2_update_0_stage_105 <= bright_gauss_blur_2_update_0_stage_104;
      bright_gauss_blur_2_update_0_stage_106 <= bright_gauss_blur_2_update_0_stage_105;
      bright_gauss_blur_2_update_0_stage_107 <= bright_gauss_blur_2_update_0_stage_106;
      bright_gauss_blur_2_update_0_stage_108 <= bright_gauss_blur_2_update_0_stage_107;
      bright_gauss_blur_2_update_0_stage_109 <= bright_gauss_blur_2_update_0_stage_108;
      bright_gauss_blur_2_update_0_stage_110 <= bright_gauss_blur_2_update_0_stage_109;
      bright_gauss_blur_2_update_0_stage_111 <= bright_gauss_blur_2_update_0_stage_110;
      bright_gauss_blur_2_update_0_stage_112 <= bright_gauss_blur_2_update_0_stage_111;
      bright_gauss_blur_2_update_0_stage_113 <= bright_gauss_blur_2_update_0_stage_112;
      bright_gauss_blur_2_update_0_stage_114 <= bright_gauss_blur_2_update_0_stage_113;
      bright_gauss_blur_2_update_0_stage_115 <= bright_gauss_blur_2_update_0_stage_114;
      bright_gauss_blur_2_update_0_stage_116 <= bright_gauss_blur_2_update_0_stage_115;
      bright_gauss_blur_2_update_0_stage_117 <= bright_gauss_blur_2_update_0_stage_116;
      bright_gauss_blur_2_update_0_stage_118 <= bright_gauss_blur_2_update_0_stage_117;
      bright_gauss_blur_2_update_0_stage_119 <= bright_gauss_blur_2_update_0_stage_118;
      bright_gauss_blur_2_update_0_stage_120 <= bright_gauss_blur_2_update_0_stage_119;
      bright_gauss_blur_2_update_0_stage_121 <= bright_gauss_blur_2_update_0_stage_120;
      bright_gauss_blur_2_update_0_stage_122 <= bright_gauss_blur_2_update_0_stage_121;
      bright_gauss_blur_2_update_0_stage_123 <= bright_gauss_blur_2_update_0_stage_122;
      bright_gauss_blur_2_update_0_stage_124 <= bright_gauss_blur_2_update_0_stage_123;
      bright_gauss_blur_2_update_0_stage_125 <= bright_gauss_blur_2_update_0_stage_124;
      bright_gauss_blur_2_update_0_stage_126 <= bright_gauss_blur_2_update_0_stage_125;
      bright_gauss_blur_2_update_0_stage_127 <= bright_gauss_blur_2_update_0_stage_126;
      bright_gauss_blur_2_update_0_stage_128 <= bright_gauss_blur_2_update_0_stage_127;
      bright_gauss_blur_2_update_0_stage_129 <= bright_gauss_blur_2_update_0_stage_128;
      bright_gauss_blur_2_update_0_stage_130 <= bright_gauss_blur_2_update_0_stage_129;
      bright_gauss_blur_2_update_0_stage_131 <= bright_gauss_blur_2_update_0_stage_130;
      bright_gauss_blur_2_update_0_stage_132 <= bright_gauss_blur_2_update_0_stage_131;
      bright_gauss_blur_2_update_0_stage_133 <= bright_gauss_blur_2_update_0_stage_132;
      bright_gauss_blur_2_update_0_stage_134 <= bright_gauss_blur_2_update_0_stage_133;
      bright_gauss_blur_2_update_0_stage_135 <= bright_gauss_blur_2_update_0_stage_134;
      bright_gauss_blur_2_update_0_stage_136 <= bright_gauss_blur_2_update_0_stage_135;
      bright_gauss_blur_2_update_0_stage_137 <= bright_gauss_blur_2_update_0_stage_136;
      bright_gauss_blur_2_update_0_stage_138 <= bright_gauss_blur_2_update_0_stage_137;
      bright_gauss_blur_2_update_0_stage_139 <= bright_gauss_blur_2_update_0_stage_138;
      bright_gauss_blur_2_update_0_stage_140 <= bright_gauss_blur_2_update_0_stage_139;
      bright_gauss_blur_2_update_0_stage_141 <= bright_gauss_blur_2_update_0_stage_140;
      bright_gauss_blur_2_update_0_stage_142 <= bright_gauss_blur_2_update_0_stage_141;
      bright_gauss_blur_2_update_0_stage_143 <= bright_gauss_blur_2_update_0_stage_142;
      bright_gauss_blur_2_update_0_stage_144 <= bright_gauss_blur_2_update_0_stage_143;
      bright_gauss_blur_2_update_0_stage_145 <= bright_gauss_blur_2_update_0_stage_144;
      bright_gauss_blur_2_update_0_stage_146 <= bright_gauss_blur_2_update_0_stage_145;
      bright_gauss_blur_2_update_0_stage_147 <= bright_gauss_blur_2_update_0_stage_146;
      bright_gauss_blur_2_update_0_stage_148 <= bright_gauss_blur_2_update_0_stage_147;
      bright_gauss_blur_2_update_0_stage_149 <= bright_gauss_blur_2_update_0_stage_148;
      bright_gauss_blur_2_update_0_stage_150 <= bright_gauss_blur_2_update_0_stage_149;
      bright_gauss_blur_2_update_0_stage_151 <= bright_gauss_blur_2_update_0_stage_150;
      bright_gauss_blur_2_update_0_stage_152 <= bright_gauss_blur_2_update_0_stage_151;
      bright_gauss_blur_2_update_0_stage_153 <= bright_gauss_blur_2_update_0_stage_152;
      bright_gauss_blur_2_update_0_stage_154 <= bright_gauss_blur_2_update_0_stage_153;
      bright_gauss_blur_2_update_0_stage_155 <= bright_gauss_blur_2_update_0_stage_154;
      bright_gauss_blur_2_update_0_stage_156 <= bright_gauss_blur_2_update_0_stage_155;
      bright_gauss_blur_2_update_0_stage_157 <= bright_gauss_blur_2_update_0_stage_156;
      bright_gauss_blur_2_update_0_stage_158 <= bright_gauss_blur_2_update_0_stage_157;
      bright_gauss_blur_2_update_0_stage_159 <= bright_gauss_blur_2_update_0_stage_158;
      bright_gauss_blur_2_update_0_stage_160 <= bright_gauss_blur_2_update_0_stage_159;
      bright_gauss_blur_2_update_0_stage_161 <= bright_gauss_blur_2_update_0_stage_160;
      bright_gauss_blur_2_update_0_stage_162 <= bright_gauss_blur_2_update_0_stage_161;
      bright_gauss_blur_2_update_0_stage_163 <= bright_gauss_blur_2_update_0_stage_162;
      bright_gauss_blur_2_update_0_stage_164 <= bright_gauss_blur_2_update_0_stage_163;
      bright_gauss_blur_2_update_0_stage_165 <= bright_gauss_blur_2_update_0_stage_164;
      bright_gauss_blur_2_update_0_stage_166 <= bright_gauss_blur_2_update_0_stage_165;
      bright_gauss_blur_2_update_0_stage_167 <= bright_gauss_blur_2_update_0_stage_166;
      bright_gauss_blur_2_update_0_stage_168 <= bright_gauss_blur_2_update_0_stage_167;
      bright_gauss_blur_2_update_0_stage_169 <= bright_gauss_blur_2_update_0_stage_168;
      bright_gauss_blur_2_update_0_stage_170 <= bright_gauss_blur_2_update_0_stage_169;
      bright_gauss_blur_2_update_0_stage_171 <= bright_gauss_blur_2_update_0_stage_170;
      bright_gauss_blur_2_update_0_stage_172 <= bright_gauss_blur_2_update_0_stage_171;
      bright_gauss_blur_2_update_0_stage_173 <= bright_gauss_blur_2_update_0_stage_172;
      bright_gauss_blur_2_update_0_stage_174 <= bright_gauss_blur_2_update_0_stage_173;
      bright_gauss_blur_2_update_0_stage_175 <= bright_gauss_blur_2_update_0_stage_174;
      bright_gauss_blur_2_update_0_stage_176 <= bright_gauss_blur_2_update_0_stage_175;
      bright_gauss_blur_2_update_0_stage_177 <= bright_gauss_blur_2_update_0_stage_176;
      bright_gauss_blur_2_update_0_stage_178 <= bright_gauss_blur_2_update_0_stage_177;
      bright_gauss_blur_2_update_0_stage_179 <= bright_gauss_blur_2_update_0_stage_178;
      bright_gauss_blur_2_update_0_stage_180 <= bright_gauss_blur_2_update_0_stage_179;
      bright_gauss_blur_2_update_0_stage_181 <= bright_gauss_blur_2_update_0_stage_180;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_41 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_42 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_41;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_43 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_42;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_44 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_43;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_45 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_44;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_46 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_45;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_47 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_46;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_48 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_47;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_49 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_48;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_50 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_49;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_51 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_50;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_52 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_51;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_53 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_52;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_54 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_53;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_55 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_54;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_56 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_55;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_57 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_56;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_58 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_57;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_59 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_58;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_60 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_59;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_61 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_60;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_62 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_61;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_63 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_62;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_64 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_63;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_65 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_64;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_66 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_65;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_67 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_66;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_68 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_67;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_69 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_68;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_70 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_69;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_71 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_70;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_72 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_71;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_73 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_72;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_74 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_73;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_75 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_74;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_76 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_75;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_77 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_76;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_78 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_77;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_79 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_78;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_80 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_79;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_81 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_80;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_82 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_81;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_83 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_82;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_84 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_83;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_85 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_84;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_86 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_85;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_87 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_86;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_88 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_87;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_89 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_88;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_90 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_89;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_91 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_90;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_92 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_91;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_93 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_92;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_94 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_93;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_95 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_94;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_96 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_95;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_97 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_96;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_98 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_97;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_99 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_98;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_100 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_99;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_101 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_100;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_102 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_101;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_103 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_102;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_104 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_103;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_105 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_104;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_106 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_105;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_107 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_106;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_108 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_107;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_109 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_108;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_110 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_109;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_111 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_110;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_112 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_111;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_113 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_112;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_114 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_113;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_115 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_114;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_116 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_115;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_117 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_116;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_118 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_117;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_119 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_118;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_120 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_119;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_121 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_120;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_122 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_121;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_123 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_122;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_124 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_123;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_125 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_124;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_126 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_125;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_127 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_126;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_128 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_127;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_129 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_128;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_130 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_129;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_131 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_130;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_132 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_131;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_133 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_132;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_134 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_133;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_135 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_134;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_136 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_135;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_137 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_136;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_138 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_137;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_139 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_138;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_140 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_139;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_141 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_140;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_142 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_141;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_143 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_142;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_144 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_143;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_145 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_144;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_146 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_145;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_147 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_146;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_148 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_147;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_149 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_148;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_150 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_149;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_151 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_150;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_152 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_151;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_153 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_152;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_154 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_153;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_155 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_154;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_156 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_155;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_157 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_156;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_158 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_157;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_159 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_158;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_160 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_159;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_161 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_160;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_162 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_161;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_163 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_162;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_164 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_163;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_165 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_164;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_166 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_165;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_167 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_166;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_168 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_167;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_169 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_168;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_170 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_169;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_171 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_170;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_172 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_171;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_173 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_172;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_174 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_173;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_175 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_174;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_176 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_175;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_177 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_176;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_178 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_177;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_179 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_178;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_180 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_179;
      bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_181 <= bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26_stage_180;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_46 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_47 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_46;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_48 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_47;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_49 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_48;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_50 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_49;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_51 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_50;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_52 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_51;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_53 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_52;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_54 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_53;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_55 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_54;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_56 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_55;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_57 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_56;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_58 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_57;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_59 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_58;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_60 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_59;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_61 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_60;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_62 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_61;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_63 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_62;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_64 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_63;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_65 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_64;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_66 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_65;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_67 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_66;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_68 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_67;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_69 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_68;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_70 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_69;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_71 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_70;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_72 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_71;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_73 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_72;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_74 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_73;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_75 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_74;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_76 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_75;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_77 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_76;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_78 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_77;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_79 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_78;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_80 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_79;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_81 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_80;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_82 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_81;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_83 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_82;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_84 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_83;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_85 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_84;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_86 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_85;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_87 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_86;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_88 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_87;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_89 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_88;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_90 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_89;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_91 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_90;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_92 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_91;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_93 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_92;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_94 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_93;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_95 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_94;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_96 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_95;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_97 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_96;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_98 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_97;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_99 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_98;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_100 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_99;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_101 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_100;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_102 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_101;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_103 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_102;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_104 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_103;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_105 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_104;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_106 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_105;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_107 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_106;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_108 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_107;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_109 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_108;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_110 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_109;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_111 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_110;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_112 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_111;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_113 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_112;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_114 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_113;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_115 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_114;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_116 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_115;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_117 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_116;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_118 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_117;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_119 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_118;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_120 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_119;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_121 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_120;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_122 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_121;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_123 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_122;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_124 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_123;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_125 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_124;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_126 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_125;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_127 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_126;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_128 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_127;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_129 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_128;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_130 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_129;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_131 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_130;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_132 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_131;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_133 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_132;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_134 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_133;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_135 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_134;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_136 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_135;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_137 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_136;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_138 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_137;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_139 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_138;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_140 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_139;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_141 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_140;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_142 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_141;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_143 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_142;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_144 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_143;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_145 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_144;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_146 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_145;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_147 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_146;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_148 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_147;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_149 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_148;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_150 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_149;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_151 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_150;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_152 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_151;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_153 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_152;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_154 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_153;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_155 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_154;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_156 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_155;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_157 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_156;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_158 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_157;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_159 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_158;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_160 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_159;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_161 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_160;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_162 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_161;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_163 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_162;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_164 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_163;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_165 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_164;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_166 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_165;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_167 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_166;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_168 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_167;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_169 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_168;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_170 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_169;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_171 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_170;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_172 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_171;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_173 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_172;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_174 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_173;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_175 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_174;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_176 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_175;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_177 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_176;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_178 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_177;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_179 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_178;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_180 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_179;
      bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_181 <= bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30_stage_180;
      bright_laplace_us_0_update_0_stage_47 <= bright_laplace_us_0_update_0;
      bright_laplace_us_0_update_0_stage_48 <= bright_laplace_us_0_update_0_stage_47;
      bright_laplace_us_0_update_0_stage_49 <= bright_laplace_us_0_update_0_stage_48;
      bright_laplace_us_0_update_0_stage_50 <= bright_laplace_us_0_update_0_stage_49;
      bright_laplace_us_0_update_0_stage_51 <= bright_laplace_us_0_update_0_stage_50;
      bright_laplace_us_0_update_0_stage_52 <= bright_laplace_us_0_update_0_stage_51;
      bright_laplace_us_0_update_0_stage_53 <= bright_laplace_us_0_update_0_stage_52;
      bright_laplace_us_0_update_0_stage_54 <= bright_laplace_us_0_update_0_stage_53;
      bright_laplace_us_0_update_0_stage_55 <= bright_laplace_us_0_update_0_stage_54;
      bright_laplace_us_0_update_0_stage_56 <= bright_laplace_us_0_update_0_stage_55;
      bright_laplace_us_0_update_0_stage_57 <= bright_laplace_us_0_update_0_stage_56;
      bright_laplace_us_0_update_0_stage_58 <= bright_laplace_us_0_update_0_stage_57;
      bright_laplace_us_0_update_0_stage_59 <= bright_laplace_us_0_update_0_stage_58;
      bright_laplace_us_0_update_0_stage_60 <= bright_laplace_us_0_update_0_stage_59;
      bright_laplace_us_0_update_0_stage_61 <= bright_laplace_us_0_update_0_stage_60;
      bright_laplace_us_0_update_0_stage_62 <= bright_laplace_us_0_update_0_stage_61;
      bright_laplace_us_0_update_0_stage_63 <= bright_laplace_us_0_update_0_stage_62;
      bright_laplace_us_0_update_0_stage_64 <= bright_laplace_us_0_update_0_stage_63;
      bright_laplace_us_0_update_0_stage_65 <= bright_laplace_us_0_update_0_stage_64;
      bright_laplace_us_0_update_0_stage_66 <= bright_laplace_us_0_update_0_stage_65;
      bright_laplace_us_0_update_0_stage_67 <= bright_laplace_us_0_update_0_stage_66;
      bright_laplace_us_0_update_0_stage_68 <= bright_laplace_us_0_update_0_stage_67;
      bright_laplace_us_0_update_0_stage_69 <= bright_laplace_us_0_update_0_stage_68;
      bright_laplace_us_0_update_0_stage_70 <= bright_laplace_us_0_update_0_stage_69;
      bright_laplace_us_0_update_0_stage_71 <= bright_laplace_us_0_update_0_stage_70;
      bright_laplace_us_0_update_0_stage_72 <= bright_laplace_us_0_update_0_stage_71;
      bright_laplace_us_0_update_0_stage_73 <= bright_laplace_us_0_update_0_stage_72;
      bright_laplace_us_0_update_0_stage_74 <= bright_laplace_us_0_update_0_stage_73;
      bright_laplace_us_0_update_0_stage_75 <= bright_laplace_us_0_update_0_stage_74;
      bright_laplace_us_0_update_0_stage_76 <= bright_laplace_us_0_update_0_stage_75;
      bright_laplace_us_0_update_0_stage_77 <= bright_laplace_us_0_update_0_stage_76;
      bright_laplace_us_0_update_0_stage_78 <= bright_laplace_us_0_update_0_stage_77;
      bright_laplace_us_0_update_0_stage_79 <= bright_laplace_us_0_update_0_stage_78;
      bright_laplace_us_0_update_0_stage_80 <= bright_laplace_us_0_update_0_stage_79;
      bright_laplace_us_0_update_0_stage_81 <= bright_laplace_us_0_update_0_stage_80;
      bright_laplace_us_0_update_0_stage_82 <= bright_laplace_us_0_update_0_stage_81;
      bright_laplace_us_0_update_0_stage_83 <= bright_laplace_us_0_update_0_stage_82;
      bright_laplace_us_0_update_0_stage_84 <= bright_laplace_us_0_update_0_stage_83;
      bright_laplace_us_0_update_0_stage_85 <= bright_laplace_us_0_update_0_stage_84;
      bright_laplace_us_0_update_0_stage_86 <= bright_laplace_us_0_update_0_stage_85;
      bright_laplace_us_0_update_0_stage_87 <= bright_laplace_us_0_update_0_stage_86;
      bright_laplace_us_0_update_0_stage_88 <= bright_laplace_us_0_update_0_stage_87;
      bright_laplace_us_0_update_0_stage_89 <= bright_laplace_us_0_update_0_stage_88;
      bright_laplace_us_0_update_0_stage_90 <= bright_laplace_us_0_update_0_stage_89;
      bright_laplace_us_0_update_0_stage_91 <= bright_laplace_us_0_update_0_stage_90;
      bright_laplace_us_0_update_0_stage_92 <= bright_laplace_us_0_update_0_stage_91;
      bright_laplace_us_0_update_0_stage_93 <= bright_laplace_us_0_update_0_stage_92;
      bright_laplace_us_0_update_0_stage_94 <= bright_laplace_us_0_update_0_stage_93;
      bright_laplace_us_0_update_0_stage_95 <= bright_laplace_us_0_update_0_stage_94;
      bright_laplace_us_0_update_0_stage_96 <= bright_laplace_us_0_update_0_stage_95;
      bright_laplace_us_0_update_0_stage_97 <= bright_laplace_us_0_update_0_stage_96;
      bright_laplace_us_0_update_0_stage_98 <= bright_laplace_us_0_update_0_stage_97;
      bright_laplace_us_0_update_0_stage_99 <= bright_laplace_us_0_update_0_stage_98;
      bright_laplace_us_0_update_0_stage_100 <= bright_laplace_us_0_update_0_stage_99;
      bright_laplace_us_0_update_0_stage_101 <= bright_laplace_us_0_update_0_stage_100;
      bright_laplace_us_0_update_0_stage_102 <= bright_laplace_us_0_update_0_stage_101;
      bright_laplace_us_0_update_0_stage_103 <= bright_laplace_us_0_update_0_stage_102;
      bright_laplace_us_0_update_0_stage_104 <= bright_laplace_us_0_update_0_stage_103;
      bright_laplace_us_0_update_0_stage_105 <= bright_laplace_us_0_update_0_stage_104;
      bright_laplace_us_0_update_0_stage_106 <= bright_laplace_us_0_update_0_stage_105;
      bright_laplace_us_0_update_0_stage_107 <= bright_laplace_us_0_update_0_stage_106;
      bright_laplace_us_0_update_0_stage_108 <= bright_laplace_us_0_update_0_stage_107;
      bright_laplace_us_0_update_0_stage_109 <= bright_laplace_us_0_update_0_stage_108;
      bright_laplace_us_0_update_0_stage_110 <= bright_laplace_us_0_update_0_stage_109;
      bright_laplace_us_0_update_0_stage_111 <= bright_laplace_us_0_update_0_stage_110;
      bright_laplace_us_0_update_0_stage_112 <= bright_laplace_us_0_update_0_stage_111;
      bright_laplace_us_0_update_0_stage_113 <= bright_laplace_us_0_update_0_stage_112;
      bright_laplace_us_0_update_0_stage_114 <= bright_laplace_us_0_update_0_stage_113;
      bright_laplace_us_0_update_0_stage_115 <= bright_laplace_us_0_update_0_stage_114;
      bright_laplace_us_0_update_0_stage_116 <= bright_laplace_us_0_update_0_stage_115;
      bright_laplace_us_0_update_0_stage_117 <= bright_laplace_us_0_update_0_stage_116;
      bright_laplace_us_0_update_0_stage_118 <= bright_laplace_us_0_update_0_stage_117;
      bright_laplace_us_0_update_0_stage_119 <= bright_laplace_us_0_update_0_stage_118;
      bright_laplace_us_0_update_0_stage_120 <= bright_laplace_us_0_update_0_stage_119;
      bright_laplace_us_0_update_0_stage_121 <= bright_laplace_us_0_update_0_stage_120;
      bright_laplace_us_0_update_0_stage_122 <= bright_laplace_us_0_update_0_stage_121;
      bright_laplace_us_0_update_0_stage_123 <= bright_laplace_us_0_update_0_stage_122;
      bright_laplace_us_0_update_0_stage_124 <= bright_laplace_us_0_update_0_stage_123;
      bright_laplace_us_0_update_0_stage_125 <= bright_laplace_us_0_update_0_stage_124;
      bright_laplace_us_0_update_0_stage_126 <= bright_laplace_us_0_update_0_stage_125;
      bright_laplace_us_0_update_0_stage_127 <= bright_laplace_us_0_update_0_stage_126;
      bright_laplace_us_0_update_0_stage_128 <= bright_laplace_us_0_update_0_stage_127;
      bright_laplace_us_0_update_0_stage_129 <= bright_laplace_us_0_update_0_stage_128;
      bright_laplace_us_0_update_0_stage_130 <= bright_laplace_us_0_update_0_stage_129;
      bright_laplace_us_0_update_0_stage_131 <= bright_laplace_us_0_update_0_stage_130;
      bright_laplace_us_0_update_0_stage_132 <= bright_laplace_us_0_update_0_stage_131;
      bright_laplace_us_0_update_0_stage_133 <= bright_laplace_us_0_update_0_stage_132;
      bright_laplace_us_0_update_0_stage_134 <= bright_laplace_us_0_update_0_stage_133;
      bright_laplace_us_0_update_0_stage_135 <= bright_laplace_us_0_update_0_stage_134;
      bright_laplace_us_0_update_0_stage_136 <= bright_laplace_us_0_update_0_stage_135;
      bright_laplace_us_0_update_0_stage_137 <= bright_laplace_us_0_update_0_stage_136;
      bright_laplace_us_0_update_0_stage_138 <= bright_laplace_us_0_update_0_stage_137;
      bright_laplace_us_0_update_0_stage_139 <= bright_laplace_us_0_update_0_stage_138;
      bright_laplace_us_0_update_0_stage_140 <= bright_laplace_us_0_update_0_stage_139;
      bright_laplace_us_0_update_0_stage_141 <= bright_laplace_us_0_update_0_stage_140;
      bright_laplace_us_0_update_0_stage_142 <= bright_laplace_us_0_update_0_stage_141;
      bright_laplace_us_0_update_0_stage_143 <= bright_laplace_us_0_update_0_stage_142;
      bright_laplace_us_0_update_0_stage_144 <= bright_laplace_us_0_update_0_stage_143;
      bright_laplace_us_0_update_0_stage_145 <= bright_laplace_us_0_update_0_stage_144;
      bright_laplace_us_0_update_0_stage_146 <= bright_laplace_us_0_update_0_stage_145;
      bright_laplace_us_0_update_0_stage_147 <= bright_laplace_us_0_update_0_stage_146;
      bright_laplace_us_0_update_0_stage_148 <= bright_laplace_us_0_update_0_stage_147;
      bright_laplace_us_0_update_0_stage_149 <= bright_laplace_us_0_update_0_stage_148;
      bright_laplace_us_0_update_0_stage_150 <= bright_laplace_us_0_update_0_stage_149;
      bright_laplace_us_0_update_0_stage_151 <= bright_laplace_us_0_update_0_stage_150;
      bright_laplace_us_0_update_0_stage_152 <= bright_laplace_us_0_update_0_stage_151;
      bright_laplace_us_0_update_0_stage_153 <= bright_laplace_us_0_update_0_stage_152;
      bright_laplace_us_0_update_0_stage_154 <= bright_laplace_us_0_update_0_stage_153;
      bright_laplace_us_0_update_0_stage_155 <= bright_laplace_us_0_update_0_stage_154;
      bright_laplace_us_0_update_0_stage_156 <= bright_laplace_us_0_update_0_stage_155;
      bright_laplace_us_0_update_0_stage_157 <= bright_laplace_us_0_update_0_stage_156;
      bright_laplace_us_0_update_0_stage_158 <= bright_laplace_us_0_update_0_stage_157;
      bright_laplace_us_0_update_0_stage_159 <= bright_laplace_us_0_update_0_stage_158;
      bright_laplace_us_0_update_0_stage_160 <= bright_laplace_us_0_update_0_stage_159;
      bright_laplace_us_0_update_0_stage_161 <= bright_laplace_us_0_update_0_stage_160;
      bright_laplace_us_0_update_0_stage_162 <= bright_laplace_us_0_update_0_stage_161;
      bright_laplace_us_0_update_0_stage_163 <= bright_laplace_us_0_update_0_stage_162;
      bright_laplace_us_0_update_0_stage_164 <= bright_laplace_us_0_update_0_stage_163;
      bright_laplace_us_0_update_0_stage_165 <= bright_laplace_us_0_update_0_stage_164;
      bright_laplace_us_0_update_0_stage_166 <= bright_laplace_us_0_update_0_stage_165;
      bright_laplace_us_0_update_0_stage_167 <= bright_laplace_us_0_update_0_stage_166;
      bright_laplace_us_0_update_0_stage_168 <= bright_laplace_us_0_update_0_stage_167;
      bright_laplace_us_0_update_0_stage_169 <= bright_laplace_us_0_update_0_stage_168;
      bright_laplace_us_0_update_0_stage_170 <= bright_laplace_us_0_update_0_stage_169;
      bright_laplace_us_0_update_0_stage_171 <= bright_laplace_us_0_update_0_stage_170;
      bright_laplace_us_0_update_0_stage_172 <= bright_laplace_us_0_update_0_stage_171;
      bright_laplace_us_0_update_0_stage_173 <= bright_laplace_us_0_update_0_stage_172;
      bright_laplace_us_0_update_0_stage_174 <= bright_laplace_us_0_update_0_stage_173;
      bright_laplace_us_0_update_0_stage_175 <= bright_laplace_us_0_update_0_stage_174;
      bright_laplace_us_0_update_0_stage_176 <= bright_laplace_us_0_update_0_stage_175;
      bright_laplace_us_0_update_0_stage_177 <= bright_laplace_us_0_update_0_stage_176;
      bright_laplace_us_0_update_0_stage_178 <= bright_laplace_us_0_update_0_stage_177;
      bright_laplace_us_0_update_0_stage_179 <= bright_laplace_us_0_update_0_stage_178;
      bright_laplace_us_0_update_0_stage_180 <= bright_laplace_us_0_update_0_stage_179;
      bright_laplace_us_0_update_0_stage_181 <= bright_laplace_us_0_update_0_stage_180;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_48 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_49 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_48;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_50 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_49;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_51 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_50;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_52 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_51;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_53 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_52;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_54 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_53;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_55 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_54;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_56 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_55;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_57 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_56;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_58 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_57;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_59 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_58;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_60 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_59;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_61 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_60;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_62 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_61;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_63 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_62;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_64 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_63;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_65 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_64;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_66 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_65;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_67 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_66;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_68 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_67;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_69 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_68;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_70 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_69;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_71 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_70;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_72 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_71;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_73 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_72;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_74 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_73;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_75 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_74;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_76 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_75;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_77 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_76;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_78 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_77;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_79 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_78;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_80 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_79;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_81 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_80;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_82 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_81;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_83 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_82;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_84 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_83;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_85 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_84;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_86 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_85;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_87 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_86;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_88 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_87;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_89 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_88;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_90 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_89;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_91 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_90;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_92 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_91;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_93 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_92;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_94 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_93;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_95 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_94;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_96 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_95;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_97 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_96;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_98 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_97;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_99 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_98;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_100 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_99;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_101 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_100;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_102 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_101;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_103 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_102;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_104 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_103;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_105 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_104;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_106 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_105;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_107 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_106;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_108 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_107;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_109 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_108;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_110 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_109;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_111 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_110;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_112 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_111;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_113 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_112;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_114 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_113;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_115 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_114;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_116 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_115;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_117 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_116;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_118 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_117;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_119 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_118;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_120 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_119;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_121 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_120;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_122 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_121;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_123 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_122;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_124 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_123;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_125 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_124;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_126 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_125;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_127 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_126;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_128 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_127;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_129 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_128;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_130 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_129;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_131 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_130;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_132 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_131;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_133 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_132;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_134 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_133;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_135 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_134;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_136 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_135;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_137 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_136;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_138 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_137;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_139 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_138;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_140 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_139;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_141 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_140;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_142 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_141;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_143 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_142;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_144 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_143;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_145 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_144;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_146 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_145;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_147 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_146;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_148 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_147;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_149 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_148;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_150 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_149;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_151 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_150;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_152 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_151;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_153 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_152;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_154 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_153;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_155 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_154;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_156 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_155;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_157 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_156;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_158 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_157;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_159 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_158;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_160 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_159;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_161 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_160;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_162 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_161;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_163 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_162;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_164 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_163;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_165 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_164;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_166 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_165;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_167 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_166;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_168 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_167;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_169 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_168;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_170 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_169;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_171 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_170;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_172 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_171;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_173 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_172;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_174 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_173;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_175 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_174;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_176 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_175;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_177 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_176;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_178 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_177;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_179 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_178;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_180 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_179;
      bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_181 <= bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31_stage_180;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_52 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_53 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_52;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_54 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_53;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_55 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_54;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_56 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_55;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_57 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_56;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_58 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_57;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_59 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_58;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_60 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_59;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_61 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_60;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_62 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_61;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_63 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_62;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_64 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_63;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_65 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_64;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_66 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_65;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_67 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_66;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_68 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_67;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_69 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_68;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_70 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_69;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_71 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_70;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_72 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_71;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_73 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_72;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_74 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_73;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_75 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_74;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_76 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_75;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_77 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_76;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_78 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_77;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_79 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_78;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_80 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_79;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_81 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_80;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_82 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_81;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_83 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_82;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_84 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_83;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_85 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_84;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_86 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_85;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_87 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_86;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_88 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_87;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_89 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_88;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_90 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_89;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_91 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_90;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_92 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_91;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_93 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_92;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_94 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_93;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_95 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_94;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_96 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_95;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_97 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_96;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_98 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_97;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_99 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_98;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_100 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_99;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_101 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_100;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_102 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_101;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_103 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_102;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_104 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_103;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_105 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_104;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_106 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_105;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_107 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_106;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_108 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_107;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_109 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_108;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_110 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_109;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_111 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_110;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_112 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_111;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_113 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_112;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_114 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_113;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_115 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_114;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_116 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_115;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_117 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_116;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_118 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_117;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_119 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_118;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_120 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_119;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_121 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_120;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_122 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_121;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_123 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_122;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_124 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_123;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_125 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_124;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_126 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_125;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_127 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_126;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_128 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_127;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_129 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_128;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_130 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_129;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_131 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_130;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_132 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_131;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_133 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_132;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_134 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_133;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_135 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_134;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_136 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_135;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_137 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_136;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_138 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_137;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_139 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_138;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_140 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_139;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_141 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_140;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_142 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_141;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_143 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_142;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_144 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_143;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_145 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_144;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_146 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_145;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_147 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_146;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_148 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_147;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_149 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_148;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_150 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_149;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_151 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_150;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_152 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_151;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_153 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_152;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_154 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_153;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_155 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_154;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_156 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_155;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_157 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_156;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_158 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_157;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_159 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_158;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_160 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_159;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_161 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_160;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_162 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_161;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_163 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_162;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_164 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_163;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_165 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_164;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_166 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_165;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_167 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_166;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_168 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_167;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_169 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_168;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_170 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_169;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_171 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_170;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_172 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_171;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_173 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_172;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_174 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_173;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_175 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_174;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_176 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_175;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_177 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_176;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_178 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_177;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_179 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_178;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_180 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_179;
      dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_181 <= dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34_stage_180;
      dark_gauss_ds_2_update_0_stage_53 <= dark_gauss_ds_2_update_0;
      dark_gauss_ds_2_update_0_stage_54 <= dark_gauss_ds_2_update_0_stage_53;
      dark_gauss_ds_2_update_0_stage_55 <= dark_gauss_ds_2_update_0_stage_54;
      dark_gauss_ds_2_update_0_stage_56 <= dark_gauss_ds_2_update_0_stage_55;
      dark_gauss_ds_2_update_0_stage_57 <= dark_gauss_ds_2_update_0_stage_56;
      dark_gauss_ds_2_update_0_stage_58 <= dark_gauss_ds_2_update_0_stage_57;
      dark_gauss_ds_2_update_0_stage_59 <= dark_gauss_ds_2_update_0_stage_58;
      dark_gauss_ds_2_update_0_stage_60 <= dark_gauss_ds_2_update_0_stage_59;
      dark_gauss_ds_2_update_0_stage_61 <= dark_gauss_ds_2_update_0_stage_60;
      dark_gauss_ds_2_update_0_stage_62 <= dark_gauss_ds_2_update_0_stage_61;
      dark_gauss_ds_2_update_0_stage_63 <= dark_gauss_ds_2_update_0_stage_62;
      dark_gauss_ds_2_update_0_stage_64 <= dark_gauss_ds_2_update_0_stage_63;
      dark_gauss_ds_2_update_0_stage_65 <= dark_gauss_ds_2_update_0_stage_64;
      dark_gauss_ds_2_update_0_stage_66 <= dark_gauss_ds_2_update_0_stage_65;
      dark_gauss_ds_2_update_0_stage_67 <= dark_gauss_ds_2_update_0_stage_66;
      dark_gauss_ds_2_update_0_stage_68 <= dark_gauss_ds_2_update_0_stage_67;
      dark_gauss_ds_2_update_0_stage_69 <= dark_gauss_ds_2_update_0_stage_68;
      dark_gauss_ds_2_update_0_stage_70 <= dark_gauss_ds_2_update_0_stage_69;
      dark_gauss_ds_2_update_0_stage_71 <= dark_gauss_ds_2_update_0_stage_70;
      dark_gauss_ds_2_update_0_stage_72 <= dark_gauss_ds_2_update_0_stage_71;
      dark_gauss_ds_2_update_0_stage_73 <= dark_gauss_ds_2_update_0_stage_72;
      dark_gauss_ds_2_update_0_stage_74 <= dark_gauss_ds_2_update_0_stage_73;
      dark_gauss_ds_2_update_0_stage_75 <= dark_gauss_ds_2_update_0_stage_74;
      dark_gauss_ds_2_update_0_stage_76 <= dark_gauss_ds_2_update_0_stage_75;
      dark_gauss_ds_2_update_0_stage_77 <= dark_gauss_ds_2_update_0_stage_76;
      dark_gauss_ds_2_update_0_stage_78 <= dark_gauss_ds_2_update_0_stage_77;
      dark_gauss_ds_2_update_0_stage_79 <= dark_gauss_ds_2_update_0_stage_78;
      dark_gauss_ds_2_update_0_stage_80 <= dark_gauss_ds_2_update_0_stage_79;
      dark_gauss_ds_2_update_0_stage_81 <= dark_gauss_ds_2_update_0_stage_80;
      dark_gauss_ds_2_update_0_stage_82 <= dark_gauss_ds_2_update_0_stage_81;
      dark_gauss_ds_2_update_0_stage_83 <= dark_gauss_ds_2_update_0_stage_82;
      dark_gauss_ds_2_update_0_stage_84 <= dark_gauss_ds_2_update_0_stage_83;
      dark_gauss_ds_2_update_0_stage_85 <= dark_gauss_ds_2_update_0_stage_84;
      dark_gauss_ds_2_update_0_stage_86 <= dark_gauss_ds_2_update_0_stage_85;
      dark_gauss_ds_2_update_0_stage_87 <= dark_gauss_ds_2_update_0_stage_86;
      dark_gauss_ds_2_update_0_stage_88 <= dark_gauss_ds_2_update_0_stage_87;
      dark_gauss_ds_2_update_0_stage_89 <= dark_gauss_ds_2_update_0_stage_88;
      dark_gauss_ds_2_update_0_stage_90 <= dark_gauss_ds_2_update_0_stage_89;
      dark_gauss_ds_2_update_0_stage_91 <= dark_gauss_ds_2_update_0_stage_90;
      dark_gauss_ds_2_update_0_stage_92 <= dark_gauss_ds_2_update_0_stage_91;
      dark_gauss_ds_2_update_0_stage_93 <= dark_gauss_ds_2_update_0_stage_92;
      dark_gauss_ds_2_update_0_stage_94 <= dark_gauss_ds_2_update_0_stage_93;
      dark_gauss_ds_2_update_0_stage_95 <= dark_gauss_ds_2_update_0_stage_94;
      dark_gauss_ds_2_update_0_stage_96 <= dark_gauss_ds_2_update_0_stage_95;
      dark_gauss_ds_2_update_0_stage_97 <= dark_gauss_ds_2_update_0_stage_96;
      dark_gauss_ds_2_update_0_stage_98 <= dark_gauss_ds_2_update_0_stage_97;
      dark_gauss_ds_2_update_0_stage_99 <= dark_gauss_ds_2_update_0_stage_98;
      dark_gauss_ds_2_update_0_stage_100 <= dark_gauss_ds_2_update_0_stage_99;
      dark_gauss_ds_2_update_0_stage_101 <= dark_gauss_ds_2_update_0_stage_100;
      dark_gauss_ds_2_update_0_stage_102 <= dark_gauss_ds_2_update_0_stage_101;
      dark_gauss_ds_2_update_0_stage_103 <= dark_gauss_ds_2_update_0_stage_102;
      dark_gauss_ds_2_update_0_stage_104 <= dark_gauss_ds_2_update_0_stage_103;
      dark_gauss_ds_2_update_0_stage_105 <= dark_gauss_ds_2_update_0_stage_104;
      dark_gauss_ds_2_update_0_stage_106 <= dark_gauss_ds_2_update_0_stage_105;
      dark_gauss_ds_2_update_0_stage_107 <= dark_gauss_ds_2_update_0_stage_106;
      dark_gauss_ds_2_update_0_stage_108 <= dark_gauss_ds_2_update_0_stage_107;
      dark_gauss_ds_2_update_0_stage_109 <= dark_gauss_ds_2_update_0_stage_108;
      dark_gauss_ds_2_update_0_stage_110 <= dark_gauss_ds_2_update_0_stage_109;
      dark_gauss_ds_2_update_0_stage_111 <= dark_gauss_ds_2_update_0_stage_110;
      dark_gauss_ds_2_update_0_stage_112 <= dark_gauss_ds_2_update_0_stage_111;
      dark_gauss_ds_2_update_0_stage_113 <= dark_gauss_ds_2_update_0_stage_112;
      dark_gauss_ds_2_update_0_stage_114 <= dark_gauss_ds_2_update_0_stage_113;
      dark_gauss_ds_2_update_0_stage_115 <= dark_gauss_ds_2_update_0_stage_114;
      dark_gauss_ds_2_update_0_stage_116 <= dark_gauss_ds_2_update_0_stage_115;
      dark_gauss_ds_2_update_0_stage_117 <= dark_gauss_ds_2_update_0_stage_116;
      dark_gauss_ds_2_update_0_stage_118 <= dark_gauss_ds_2_update_0_stage_117;
      dark_gauss_ds_2_update_0_stage_119 <= dark_gauss_ds_2_update_0_stage_118;
      dark_gauss_ds_2_update_0_stage_120 <= dark_gauss_ds_2_update_0_stage_119;
      dark_gauss_ds_2_update_0_stage_121 <= dark_gauss_ds_2_update_0_stage_120;
      dark_gauss_ds_2_update_0_stage_122 <= dark_gauss_ds_2_update_0_stage_121;
      dark_gauss_ds_2_update_0_stage_123 <= dark_gauss_ds_2_update_0_stage_122;
      dark_gauss_ds_2_update_0_stage_124 <= dark_gauss_ds_2_update_0_stage_123;
      dark_gauss_ds_2_update_0_stage_125 <= dark_gauss_ds_2_update_0_stage_124;
      dark_gauss_ds_2_update_0_stage_126 <= dark_gauss_ds_2_update_0_stage_125;
      dark_gauss_ds_2_update_0_stage_127 <= dark_gauss_ds_2_update_0_stage_126;
      dark_gauss_ds_2_update_0_stage_128 <= dark_gauss_ds_2_update_0_stage_127;
      dark_gauss_ds_2_update_0_stage_129 <= dark_gauss_ds_2_update_0_stage_128;
      dark_gauss_ds_2_update_0_stage_130 <= dark_gauss_ds_2_update_0_stage_129;
      dark_gauss_ds_2_update_0_stage_131 <= dark_gauss_ds_2_update_0_stage_130;
      dark_gauss_ds_2_update_0_stage_132 <= dark_gauss_ds_2_update_0_stage_131;
      dark_gauss_ds_2_update_0_stage_133 <= dark_gauss_ds_2_update_0_stage_132;
      dark_gauss_ds_2_update_0_stage_134 <= dark_gauss_ds_2_update_0_stage_133;
      dark_gauss_ds_2_update_0_stage_135 <= dark_gauss_ds_2_update_0_stage_134;
      dark_gauss_ds_2_update_0_stage_136 <= dark_gauss_ds_2_update_0_stage_135;
      dark_gauss_ds_2_update_0_stage_137 <= dark_gauss_ds_2_update_0_stage_136;
      dark_gauss_ds_2_update_0_stage_138 <= dark_gauss_ds_2_update_0_stage_137;
      dark_gauss_ds_2_update_0_stage_139 <= dark_gauss_ds_2_update_0_stage_138;
      dark_gauss_ds_2_update_0_stage_140 <= dark_gauss_ds_2_update_0_stage_139;
      dark_gauss_ds_2_update_0_stage_141 <= dark_gauss_ds_2_update_0_stage_140;
      dark_gauss_ds_2_update_0_stage_142 <= dark_gauss_ds_2_update_0_stage_141;
      dark_gauss_ds_2_update_0_stage_143 <= dark_gauss_ds_2_update_0_stage_142;
      dark_gauss_ds_2_update_0_stage_144 <= dark_gauss_ds_2_update_0_stage_143;
      dark_gauss_ds_2_update_0_stage_145 <= dark_gauss_ds_2_update_0_stage_144;
      dark_gauss_ds_2_update_0_stage_146 <= dark_gauss_ds_2_update_0_stage_145;
      dark_gauss_ds_2_update_0_stage_147 <= dark_gauss_ds_2_update_0_stage_146;
      dark_gauss_ds_2_update_0_stage_148 <= dark_gauss_ds_2_update_0_stage_147;
      dark_gauss_ds_2_update_0_stage_149 <= dark_gauss_ds_2_update_0_stage_148;
      dark_gauss_ds_2_update_0_stage_150 <= dark_gauss_ds_2_update_0_stage_149;
      dark_gauss_ds_2_update_0_stage_151 <= dark_gauss_ds_2_update_0_stage_150;
      dark_gauss_ds_2_update_0_stage_152 <= dark_gauss_ds_2_update_0_stage_151;
      dark_gauss_ds_2_update_0_stage_153 <= dark_gauss_ds_2_update_0_stage_152;
      dark_gauss_ds_2_update_0_stage_154 <= dark_gauss_ds_2_update_0_stage_153;
      dark_gauss_ds_2_update_0_stage_155 <= dark_gauss_ds_2_update_0_stage_154;
      dark_gauss_ds_2_update_0_stage_156 <= dark_gauss_ds_2_update_0_stage_155;
      dark_gauss_ds_2_update_0_stage_157 <= dark_gauss_ds_2_update_0_stage_156;
      dark_gauss_ds_2_update_0_stage_158 <= dark_gauss_ds_2_update_0_stage_157;
      dark_gauss_ds_2_update_0_stage_159 <= dark_gauss_ds_2_update_0_stage_158;
      dark_gauss_ds_2_update_0_stage_160 <= dark_gauss_ds_2_update_0_stage_159;
      dark_gauss_ds_2_update_0_stage_161 <= dark_gauss_ds_2_update_0_stage_160;
      dark_gauss_ds_2_update_0_stage_162 <= dark_gauss_ds_2_update_0_stage_161;
      dark_gauss_ds_2_update_0_stage_163 <= dark_gauss_ds_2_update_0_stage_162;
      dark_gauss_ds_2_update_0_stage_164 <= dark_gauss_ds_2_update_0_stage_163;
      dark_gauss_ds_2_update_0_stage_165 <= dark_gauss_ds_2_update_0_stage_164;
      dark_gauss_ds_2_update_0_stage_166 <= dark_gauss_ds_2_update_0_stage_165;
      dark_gauss_ds_2_update_0_stage_167 <= dark_gauss_ds_2_update_0_stage_166;
      dark_gauss_ds_2_update_0_stage_168 <= dark_gauss_ds_2_update_0_stage_167;
      dark_gauss_ds_2_update_0_stage_169 <= dark_gauss_ds_2_update_0_stage_168;
      dark_gauss_ds_2_update_0_stage_170 <= dark_gauss_ds_2_update_0_stage_169;
      dark_gauss_ds_2_update_0_stage_171 <= dark_gauss_ds_2_update_0_stage_170;
      dark_gauss_ds_2_update_0_stage_172 <= dark_gauss_ds_2_update_0_stage_171;
      dark_gauss_ds_2_update_0_stage_173 <= dark_gauss_ds_2_update_0_stage_172;
      dark_gauss_ds_2_update_0_stage_174 <= dark_gauss_ds_2_update_0_stage_173;
      dark_gauss_ds_2_update_0_stage_175 <= dark_gauss_ds_2_update_0_stage_174;
      dark_gauss_ds_2_update_0_stage_176 <= dark_gauss_ds_2_update_0_stage_175;
      dark_gauss_ds_2_update_0_stage_177 <= dark_gauss_ds_2_update_0_stage_176;
      dark_gauss_ds_2_update_0_stage_178 <= dark_gauss_ds_2_update_0_stage_177;
      dark_gauss_ds_2_update_0_stage_179 <= dark_gauss_ds_2_update_0_stage_178;
      dark_gauss_ds_2_update_0_stage_180 <= dark_gauss_ds_2_update_0_stage_179;
      dark_gauss_ds_2_update_0_stage_181 <= dark_gauss_ds_2_update_0_stage_180;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_54 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_55 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_54;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_56 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_55;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_57 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_56;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_58 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_57;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_59 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_58;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_60 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_59;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_61 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_60;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_62 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_61;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_63 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_62;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_64 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_63;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_65 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_64;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_66 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_65;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_67 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_66;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_68 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_67;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_69 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_68;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_70 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_69;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_71 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_70;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_72 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_71;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_73 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_72;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_74 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_73;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_75 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_74;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_76 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_75;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_77 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_76;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_78 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_77;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_79 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_78;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_80 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_79;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_81 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_80;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_82 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_81;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_83 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_82;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_84 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_83;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_85 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_84;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_86 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_85;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_87 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_86;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_88 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_87;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_89 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_88;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_90 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_89;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_91 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_90;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_92 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_91;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_93 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_92;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_94 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_93;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_95 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_94;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_96 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_95;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_97 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_96;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_98 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_97;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_99 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_98;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_100 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_99;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_101 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_100;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_102 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_101;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_103 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_102;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_104 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_103;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_105 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_104;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_106 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_105;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_107 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_106;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_108 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_107;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_109 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_108;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_110 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_109;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_111 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_110;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_112 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_111;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_113 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_112;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_114 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_113;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_115 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_114;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_116 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_115;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_117 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_116;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_118 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_117;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_119 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_118;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_120 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_119;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_121 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_120;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_122 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_121;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_123 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_122;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_124 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_123;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_125 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_124;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_126 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_125;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_127 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_126;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_128 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_127;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_129 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_128;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_130 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_129;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_131 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_130;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_132 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_131;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_133 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_132;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_134 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_133;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_135 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_134;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_136 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_135;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_137 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_136;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_138 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_137;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_139 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_138;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_140 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_139;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_141 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_140;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_142 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_141;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_143 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_142;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_144 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_143;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_145 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_144;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_146 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_145;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_147 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_146;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_148 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_147;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_149 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_148;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_150 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_149;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_151 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_150;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_152 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_151;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_153 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_152;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_154 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_153;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_155 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_154;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_156 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_155;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_157 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_156;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_158 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_157;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_159 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_158;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_160 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_159;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_161 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_160;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_162 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_161;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_163 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_162;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_164 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_163;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_165 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_164;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_166 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_165;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_167 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_166;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_168 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_167;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_169 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_168;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_170 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_169;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_171 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_170;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_172 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_171;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_173 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_172;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_174 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_173;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_175 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_174;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_176 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_175;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_177 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_176;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_178 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_177;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_179 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_178;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_180 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_179;
      dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_181 <= dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35_stage_180;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_107 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_108 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_107;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_109 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_108;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_110 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_109;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_111 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_110;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_112 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_111;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_113 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_112;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_114 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_113;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_115 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_114;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_116 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_115;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_117 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_116;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_118 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_117;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_119 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_118;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_120 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_119;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_121 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_120;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_122 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_121;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_123 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_122;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_124 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_123;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_125 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_124;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_126 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_125;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_127 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_126;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_128 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_127;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_129 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_128;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_130 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_129;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_131 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_130;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_132 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_131;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_133 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_132;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_134 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_133;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_135 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_134;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_136 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_135;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_137 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_136;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_138 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_137;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_139 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_138;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_140 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_139;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_141 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_140;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_142 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_141;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_143 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_142;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_144 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_143;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_145 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_144;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_146 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_145;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_147 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_146;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_148 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_147;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_149 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_148;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_150 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_149;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_151 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_150;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_152 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_151;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_153 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_152;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_154 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_153;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_155 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_154;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_156 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_155;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_157 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_156;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_158 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_157;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_159 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_158;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_160 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_159;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_161 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_160;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_162 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_161;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_163 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_162;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_164 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_163;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_165 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_164;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_166 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_165;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_167 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_166;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_168 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_167;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_169 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_168;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_170 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_169;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_171 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_170;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_172 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_171;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_173 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_172;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_174 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_173;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_175 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_174;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_176 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_175;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_177 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_176;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_178 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_177;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_179 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_178;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_180 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_179;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_181 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72_stage_180;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_55 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_56 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_55;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_57 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_56;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_58 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_57;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_59 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_58;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_60 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_59;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_61 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_60;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_62 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_61;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_63 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_62;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_64 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_63;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_65 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_64;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_66 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_65;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_67 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_66;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_68 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_67;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_69 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_68;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_70 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_69;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_71 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_70;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_72 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_71;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_73 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_72;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_74 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_73;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_75 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_74;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_76 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_75;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_77 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_76;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_78 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_77;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_79 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_78;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_80 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_79;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_81 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_80;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_82 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_81;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_83 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_82;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_84 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_83;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_85 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_84;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_86 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_85;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_87 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_86;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_88 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_87;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_89 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_88;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_90 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_89;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_91 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_90;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_92 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_91;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_93 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_92;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_94 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_93;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_95 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_94;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_96 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_95;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_97 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_96;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_98 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_97;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_99 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_98;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_100 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_99;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_101 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_100;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_102 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_101;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_103 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_102;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_104 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_103;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_105 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_104;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_106 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_105;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_107 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_106;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_108 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_107;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_109 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_108;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_110 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_109;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_111 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_110;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_112 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_111;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_113 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_112;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_114 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_113;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_115 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_114;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_116 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_115;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_117 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_116;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_118 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_117;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_119 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_118;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_120 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_119;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_121 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_120;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_122 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_121;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_123 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_122;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_124 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_123;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_125 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_124;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_126 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_125;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_127 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_126;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_128 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_127;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_129 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_128;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_130 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_129;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_131 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_130;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_132 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_131;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_133 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_132;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_134 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_133;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_135 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_134;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_136 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_135;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_137 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_136;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_138 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_137;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_139 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_138;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_140 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_139;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_141 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_140;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_142 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_141;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_143 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_142;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_144 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_143;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_145 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_144;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_146 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_145;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_147 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_146;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_148 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_147;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_149 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_148;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_150 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_149;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_151 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_150;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_152 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_151;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_153 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_152;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_154 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_153;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_155 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_154;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_156 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_155;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_157 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_156;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_158 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_157;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_159 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_158;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_160 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_159;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_161 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_160;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_162 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_161;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_163 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_162;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_164 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_163;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_165 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_164;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_166 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_165;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_167 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_166;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_168 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_167;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_169 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_168;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_170 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_169;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_171 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_170;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_172 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_171;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_173 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_172;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_174 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_173;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_175 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_174;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_176 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_175;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_177 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_176;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_178 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_177;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_179 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_178;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_180 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_179;
      bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_181 <= bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36_stage_180;
      bright_gauss_blur_3_update_0_stage_56 <= bright_gauss_blur_3_update_0;
      bright_gauss_blur_3_update_0_stage_57 <= bright_gauss_blur_3_update_0_stage_56;
      bright_gauss_blur_3_update_0_stage_58 <= bright_gauss_blur_3_update_0_stage_57;
      bright_gauss_blur_3_update_0_stage_59 <= bright_gauss_blur_3_update_0_stage_58;
      bright_gauss_blur_3_update_0_stage_60 <= bright_gauss_blur_3_update_0_stage_59;
      bright_gauss_blur_3_update_0_stage_61 <= bright_gauss_blur_3_update_0_stage_60;
      bright_gauss_blur_3_update_0_stage_62 <= bright_gauss_blur_3_update_0_stage_61;
      bright_gauss_blur_3_update_0_stage_63 <= bright_gauss_blur_3_update_0_stage_62;
      bright_gauss_blur_3_update_0_stage_64 <= bright_gauss_blur_3_update_0_stage_63;
      bright_gauss_blur_3_update_0_stage_65 <= bright_gauss_blur_3_update_0_stage_64;
      bright_gauss_blur_3_update_0_stage_66 <= bright_gauss_blur_3_update_0_stage_65;
      bright_gauss_blur_3_update_0_stage_67 <= bright_gauss_blur_3_update_0_stage_66;
      bright_gauss_blur_3_update_0_stage_68 <= bright_gauss_blur_3_update_0_stage_67;
      bright_gauss_blur_3_update_0_stage_69 <= bright_gauss_blur_3_update_0_stage_68;
      bright_gauss_blur_3_update_0_stage_70 <= bright_gauss_blur_3_update_0_stage_69;
      bright_gauss_blur_3_update_0_stage_71 <= bright_gauss_blur_3_update_0_stage_70;
      bright_gauss_blur_3_update_0_stage_72 <= bright_gauss_blur_3_update_0_stage_71;
      bright_gauss_blur_3_update_0_stage_73 <= bright_gauss_blur_3_update_0_stage_72;
      bright_gauss_blur_3_update_0_stage_74 <= bright_gauss_blur_3_update_0_stage_73;
      bright_gauss_blur_3_update_0_stage_75 <= bright_gauss_blur_3_update_0_stage_74;
      bright_gauss_blur_3_update_0_stage_76 <= bright_gauss_blur_3_update_0_stage_75;
      bright_gauss_blur_3_update_0_stage_77 <= bright_gauss_blur_3_update_0_stage_76;
      bright_gauss_blur_3_update_0_stage_78 <= bright_gauss_blur_3_update_0_stage_77;
      bright_gauss_blur_3_update_0_stage_79 <= bright_gauss_blur_3_update_0_stage_78;
      bright_gauss_blur_3_update_0_stage_80 <= bright_gauss_blur_3_update_0_stage_79;
      bright_gauss_blur_3_update_0_stage_81 <= bright_gauss_blur_3_update_0_stage_80;
      bright_gauss_blur_3_update_0_stage_82 <= bright_gauss_blur_3_update_0_stage_81;
      bright_gauss_blur_3_update_0_stage_83 <= bright_gauss_blur_3_update_0_stage_82;
      bright_gauss_blur_3_update_0_stage_84 <= bright_gauss_blur_3_update_0_stage_83;
      bright_gauss_blur_3_update_0_stage_85 <= bright_gauss_blur_3_update_0_stage_84;
      bright_gauss_blur_3_update_0_stage_86 <= bright_gauss_blur_3_update_0_stage_85;
      bright_gauss_blur_3_update_0_stage_87 <= bright_gauss_blur_3_update_0_stage_86;
      bright_gauss_blur_3_update_0_stage_88 <= bright_gauss_blur_3_update_0_stage_87;
      bright_gauss_blur_3_update_0_stage_89 <= bright_gauss_blur_3_update_0_stage_88;
      bright_gauss_blur_3_update_0_stage_90 <= bright_gauss_blur_3_update_0_stage_89;
      bright_gauss_blur_3_update_0_stage_91 <= bright_gauss_blur_3_update_0_stage_90;
      bright_gauss_blur_3_update_0_stage_92 <= bright_gauss_blur_3_update_0_stage_91;
      bright_gauss_blur_3_update_0_stage_93 <= bright_gauss_blur_3_update_0_stage_92;
      bright_gauss_blur_3_update_0_stage_94 <= bright_gauss_blur_3_update_0_stage_93;
      bright_gauss_blur_3_update_0_stage_95 <= bright_gauss_blur_3_update_0_stage_94;
      bright_gauss_blur_3_update_0_stage_96 <= bright_gauss_blur_3_update_0_stage_95;
      bright_gauss_blur_3_update_0_stage_97 <= bright_gauss_blur_3_update_0_stage_96;
      bright_gauss_blur_3_update_0_stage_98 <= bright_gauss_blur_3_update_0_stage_97;
      bright_gauss_blur_3_update_0_stage_99 <= bright_gauss_blur_3_update_0_stage_98;
      bright_gauss_blur_3_update_0_stage_100 <= bright_gauss_blur_3_update_0_stage_99;
      bright_gauss_blur_3_update_0_stage_101 <= bright_gauss_blur_3_update_0_stage_100;
      bright_gauss_blur_3_update_0_stage_102 <= bright_gauss_blur_3_update_0_stage_101;
      bright_gauss_blur_3_update_0_stage_103 <= bright_gauss_blur_3_update_0_stage_102;
      bright_gauss_blur_3_update_0_stage_104 <= bright_gauss_blur_3_update_0_stage_103;
      bright_gauss_blur_3_update_0_stage_105 <= bright_gauss_blur_3_update_0_stage_104;
      bright_gauss_blur_3_update_0_stage_106 <= bright_gauss_blur_3_update_0_stage_105;
      bright_gauss_blur_3_update_0_stage_107 <= bright_gauss_blur_3_update_0_stage_106;
      bright_gauss_blur_3_update_0_stage_108 <= bright_gauss_blur_3_update_0_stage_107;
      bright_gauss_blur_3_update_0_stage_109 <= bright_gauss_blur_3_update_0_stage_108;
      bright_gauss_blur_3_update_0_stage_110 <= bright_gauss_blur_3_update_0_stage_109;
      bright_gauss_blur_3_update_0_stage_111 <= bright_gauss_blur_3_update_0_stage_110;
      bright_gauss_blur_3_update_0_stage_112 <= bright_gauss_blur_3_update_0_stage_111;
      bright_gauss_blur_3_update_0_stage_113 <= bright_gauss_blur_3_update_0_stage_112;
      bright_gauss_blur_3_update_0_stage_114 <= bright_gauss_blur_3_update_0_stage_113;
      bright_gauss_blur_3_update_0_stage_115 <= bright_gauss_blur_3_update_0_stage_114;
      bright_gauss_blur_3_update_0_stage_116 <= bright_gauss_blur_3_update_0_stage_115;
      bright_gauss_blur_3_update_0_stage_117 <= bright_gauss_blur_3_update_0_stage_116;
      bright_gauss_blur_3_update_0_stage_118 <= bright_gauss_blur_3_update_0_stage_117;
      bright_gauss_blur_3_update_0_stage_119 <= bright_gauss_blur_3_update_0_stage_118;
      bright_gauss_blur_3_update_0_stage_120 <= bright_gauss_blur_3_update_0_stage_119;
      bright_gauss_blur_3_update_0_stage_121 <= bright_gauss_blur_3_update_0_stage_120;
      bright_gauss_blur_3_update_0_stage_122 <= bright_gauss_blur_3_update_0_stage_121;
      bright_gauss_blur_3_update_0_stage_123 <= bright_gauss_blur_3_update_0_stage_122;
      bright_gauss_blur_3_update_0_stage_124 <= bright_gauss_blur_3_update_0_stage_123;
      bright_gauss_blur_3_update_0_stage_125 <= bright_gauss_blur_3_update_0_stage_124;
      bright_gauss_blur_3_update_0_stage_126 <= bright_gauss_blur_3_update_0_stage_125;
      bright_gauss_blur_3_update_0_stage_127 <= bright_gauss_blur_3_update_0_stage_126;
      bright_gauss_blur_3_update_0_stage_128 <= bright_gauss_blur_3_update_0_stage_127;
      bright_gauss_blur_3_update_0_stage_129 <= bright_gauss_blur_3_update_0_stage_128;
      bright_gauss_blur_3_update_0_stage_130 <= bright_gauss_blur_3_update_0_stage_129;
      bright_gauss_blur_3_update_0_stage_131 <= bright_gauss_blur_3_update_0_stage_130;
      bright_gauss_blur_3_update_0_stage_132 <= bright_gauss_blur_3_update_0_stage_131;
      bright_gauss_blur_3_update_0_stage_133 <= bright_gauss_blur_3_update_0_stage_132;
      bright_gauss_blur_3_update_0_stage_134 <= bright_gauss_blur_3_update_0_stage_133;
      bright_gauss_blur_3_update_0_stage_135 <= bright_gauss_blur_3_update_0_stage_134;
      bright_gauss_blur_3_update_0_stage_136 <= bright_gauss_blur_3_update_0_stage_135;
      bright_gauss_blur_3_update_0_stage_137 <= bright_gauss_blur_3_update_0_stage_136;
      bright_gauss_blur_3_update_0_stage_138 <= bright_gauss_blur_3_update_0_stage_137;
      bright_gauss_blur_3_update_0_stage_139 <= bright_gauss_blur_3_update_0_stage_138;
      bright_gauss_blur_3_update_0_stage_140 <= bright_gauss_blur_3_update_0_stage_139;
      bright_gauss_blur_3_update_0_stage_141 <= bright_gauss_blur_3_update_0_stage_140;
      bright_gauss_blur_3_update_0_stage_142 <= bright_gauss_blur_3_update_0_stage_141;
      bright_gauss_blur_3_update_0_stage_143 <= bright_gauss_blur_3_update_0_stage_142;
      bright_gauss_blur_3_update_0_stage_144 <= bright_gauss_blur_3_update_0_stage_143;
      bright_gauss_blur_3_update_0_stage_145 <= bright_gauss_blur_3_update_0_stage_144;
      bright_gauss_blur_3_update_0_stage_146 <= bright_gauss_blur_3_update_0_stage_145;
      bright_gauss_blur_3_update_0_stage_147 <= bright_gauss_blur_3_update_0_stage_146;
      bright_gauss_blur_3_update_0_stage_148 <= bright_gauss_blur_3_update_0_stage_147;
      bright_gauss_blur_3_update_0_stage_149 <= bright_gauss_blur_3_update_0_stage_148;
      bright_gauss_blur_3_update_0_stage_150 <= bright_gauss_blur_3_update_0_stage_149;
      bright_gauss_blur_3_update_0_stage_151 <= bright_gauss_blur_3_update_0_stage_150;
      bright_gauss_blur_3_update_0_stage_152 <= bright_gauss_blur_3_update_0_stage_151;
      bright_gauss_blur_3_update_0_stage_153 <= bright_gauss_blur_3_update_0_stage_152;
      bright_gauss_blur_3_update_0_stage_154 <= bright_gauss_blur_3_update_0_stage_153;
      bright_gauss_blur_3_update_0_stage_155 <= bright_gauss_blur_3_update_0_stage_154;
      bright_gauss_blur_3_update_0_stage_156 <= bright_gauss_blur_3_update_0_stage_155;
      bright_gauss_blur_3_update_0_stage_157 <= bright_gauss_blur_3_update_0_stage_156;
      bright_gauss_blur_3_update_0_stage_158 <= bright_gauss_blur_3_update_0_stage_157;
      bright_gauss_blur_3_update_0_stage_159 <= bright_gauss_blur_3_update_0_stage_158;
      bright_gauss_blur_3_update_0_stage_160 <= bright_gauss_blur_3_update_0_stage_159;
      bright_gauss_blur_3_update_0_stage_161 <= bright_gauss_blur_3_update_0_stage_160;
      bright_gauss_blur_3_update_0_stage_162 <= bright_gauss_blur_3_update_0_stage_161;
      bright_gauss_blur_3_update_0_stage_163 <= bright_gauss_blur_3_update_0_stage_162;
      bright_gauss_blur_3_update_0_stage_164 <= bright_gauss_blur_3_update_0_stage_163;
      bright_gauss_blur_3_update_0_stage_165 <= bright_gauss_blur_3_update_0_stage_164;
      bright_gauss_blur_3_update_0_stage_166 <= bright_gauss_blur_3_update_0_stage_165;
      bright_gauss_blur_3_update_0_stage_167 <= bright_gauss_blur_3_update_0_stage_166;
      bright_gauss_blur_3_update_0_stage_168 <= bright_gauss_blur_3_update_0_stage_167;
      bright_gauss_blur_3_update_0_stage_169 <= bright_gauss_blur_3_update_0_stage_168;
      bright_gauss_blur_3_update_0_stage_170 <= bright_gauss_blur_3_update_0_stage_169;
      bright_gauss_blur_3_update_0_stage_171 <= bright_gauss_blur_3_update_0_stage_170;
      bright_gauss_blur_3_update_0_stage_172 <= bright_gauss_blur_3_update_0_stage_171;
      bright_gauss_blur_3_update_0_stage_173 <= bright_gauss_blur_3_update_0_stage_172;
      bright_gauss_blur_3_update_0_stage_174 <= bright_gauss_blur_3_update_0_stage_173;
      bright_gauss_blur_3_update_0_stage_175 <= bright_gauss_blur_3_update_0_stage_174;
      bright_gauss_blur_3_update_0_stage_176 <= bright_gauss_blur_3_update_0_stage_175;
      bright_gauss_blur_3_update_0_stage_177 <= bright_gauss_blur_3_update_0_stage_176;
      bright_gauss_blur_3_update_0_stage_178 <= bright_gauss_blur_3_update_0_stage_177;
      bright_gauss_blur_3_update_0_stage_179 <= bright_gauss_blur_3_update_0_stage_178;
      bright_gauss_blur_3_update_0_stage_180 <= bright_gauss_blur_3_update_0_stage_179;
      bright_gauss_blur_3_update_0_stage_181 <= bright_gauss_blur_3_update_0_stage_180;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_57 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_58 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_57;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_59 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_58;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_60 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_59;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_61 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_60;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_62 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_61;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_63 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_62;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_64 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_63;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_65 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_64;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_66 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_65;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_67 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_66;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_68 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_67;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_69 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_68;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_70 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_69;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_71 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_70;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_72 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_71;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_73 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_72;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_74 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_73;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_75 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_74;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_76 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_75;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_77 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_76;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_78 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_77;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_79 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_78;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_80 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_79;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_81 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_80;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_82 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_81;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_83 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_82;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_84 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_83;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_85 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_84;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_86 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_85;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_87 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_86;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_88 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_87;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_89 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_88;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_90 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_89;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_91 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_90;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_92 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_91;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_93 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_92;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_94 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_93;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_95 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_94;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_96 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_95;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_97 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_96;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_98 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_97;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_99 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_98;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_100 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_99;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_101 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_100;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_102 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_101;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_103 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_102;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_104 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_103;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_105 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_104;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_106 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_105;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_107 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_106;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_108 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_107;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_109 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_108;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_110 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_109;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_111 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_110;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_112 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_111;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_113 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_112;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_114 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_113;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_115 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_114;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_116 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_115;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_117 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_116;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_118 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_117;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_119 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_118;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_120 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_119;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_121 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_120;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_122 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_121;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_123 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_122;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_124 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_123;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_125 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_124;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_126 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_125;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_127 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_126;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_128 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_127;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_129 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_128;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_130 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_129;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_131 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_130;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_132 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_131;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_133 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_132;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_134 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_133;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_135 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_134;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_136 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_135;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_137 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_136;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_138 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_137;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_139 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_138;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_140 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_139;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_141 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_140;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_142 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_141;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_143 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_142;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_144 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_143;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_145 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_144;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_146 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_145;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_147 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_146;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_148 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_147;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_149 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_148;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_150 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_149;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_151 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_150;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_152 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_151;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_153 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_152;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_154 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_153;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_155 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_154;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_156 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_155;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_157 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_156;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_158 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_157;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_159 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_158;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_160 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_159;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_161 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_160;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_162 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_161;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_163 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_162;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_164 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_163;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_165 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_164;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_166 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_165;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_167 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_166;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_168 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_167;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_169 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_168;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_170 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_169;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_171 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_170;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_172 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_171;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_173 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_172;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_174 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_173;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_175 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_174;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_176 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_175;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_177 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_176;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_178 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_177;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_179 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_178;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_180 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_179;
      bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_181 <= bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37_stage_180;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_68 <= dark_weights_dark_weights_normed_update_0_read_read_45;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_69 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_68;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_70 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_69;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_71 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_70;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_72 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_71;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_73 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_72;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_74 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_73;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_75 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_74;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_76 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_75;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_77 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_76;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_78 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_77;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_79 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_78;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_80 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_79;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_81 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_80;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_82 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_81;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_83 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_82;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_84 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_83;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_85 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_84;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_86 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_85;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_87 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_86;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_88 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_87;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_89 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_88;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_90 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_89;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_91 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_90;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_92 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_91;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_93 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_92;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_94 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_93;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_95 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_94;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_96 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_95;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_97 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_96;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_98 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_97;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_99 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_98;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_100 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_99;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_101 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_100;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_102 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_101;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_103 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_102;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_104 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_103;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_105 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_104;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_106 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_105;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_107 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_106;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_108 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_107;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_109 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_108;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_110 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_109;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_111 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_110;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_112 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_111;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_113 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_112;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_114 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_113;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_115 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_114;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_116 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_115;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_117 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_116;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_118 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_117;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_119 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_118;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_120 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_119;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_121 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_120;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_122 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_121;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_123 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_122;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_124 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_123;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_125 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_124;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_126 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_125;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_127 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_126;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_128 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_127;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_129 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_128;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_130 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_129;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_131 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_130;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_132 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_131;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_133 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_132;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_134 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_133;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_135 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_134;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_136 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_135;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_137 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_136;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_138 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_137;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_139 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_138;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_140 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_139;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_141 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_140;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_142 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_141;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_143 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_142;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_144 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_143;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_145 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_144;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_146 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_145;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_147 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_146;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_148 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_147;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_149 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_148;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_150 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_149;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_151 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_150;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_152 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_151;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_153 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_152;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_154 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_153;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_155 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_154;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_156 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_155;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_157 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_156;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_158 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_157;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_159 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_158;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_160 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_159;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_161 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_160;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_162 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_161;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_163 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_162;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_164 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_163;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_165 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_164;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_166 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_165;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_167 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_166;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_168 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_167;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_169 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_168;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_170 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_169;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_171 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_170;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_172 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_171;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_173 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_172;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_174 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_173;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_175 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_174;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_176 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_175;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_177 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_176;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_178 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_177;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_179 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_178;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_180 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_179;
      dark_weights_dark_weights_normed_update_0_read_read_45_stage_181 <= dark_weights_dark_weights_normed_update_0_read_read_45_stage_180;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_71 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_72 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_71;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_73 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_72;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_74 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_73;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_75 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_74;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_76 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_75;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_77 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_76;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_78 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_77;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_79 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_78;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_80 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_79;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_81 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_80;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_82 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_81;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_83 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_82;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_84 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_83;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_85 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_84;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_86 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_85;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_87 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_86;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_88 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_87;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_89 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_88;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_90 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_89;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_91 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_90;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_92 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_91;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_93 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_92;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_94 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_93;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_95 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_94;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_96 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_95;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_97 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_96;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_98 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_97;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_99 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_98;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_100 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_99;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_101 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_100;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_102 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_101;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_103 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_102;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_104 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_103;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_105 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_104;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_106 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_105;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_107 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_106;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_108 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_107;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_109 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_108;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_110 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_109;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_111 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_110;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_112 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_111;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_113 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_112;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_114 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_113;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_115 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_114;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_116 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_115;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_117 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_116;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_118 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_117;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_119 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_118;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_120 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_119;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_121 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_120;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_122 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_121;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_123 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_122;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_124 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_123;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_125 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_124;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_126 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_125;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_127 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_126;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_128 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_127;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_129 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_128;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_130 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_129;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_131 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_130;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_132 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_131;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_133 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_132;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_134 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_133;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_135 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_134;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_136 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_135;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_137 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_136;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_138 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_137;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_139 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_138;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_140 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_139;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_141 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_140;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_142 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_141;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_143 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_142;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_144 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_143;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_145 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_144;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_146 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_145;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_147 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_146;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_148 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_147;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_149 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_148;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_150 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_149;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_151 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_150;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_152 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_151;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_153 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_152;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_154 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_153;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_155 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_154;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_156 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_155;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_157 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_156;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_158 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_157;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_159 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_158;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_160 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_159;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_161 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_160;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_162 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_161;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_163 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_162;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_164 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_163;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_165 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_164;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_166 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_165;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_167 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_166;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_168 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_167;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_169 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_168;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_170 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_169;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_171 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_170;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_172 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_171;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_173 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_172;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_174 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_173;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_175 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_174;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_176 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_175;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_177 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_176;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_178 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_177;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_179 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_178;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_180 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_179;
      dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_181 <= dark_weights_normed_dark_weights_normed_update_0_write_write_47_stage_180;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_76 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_77 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_76;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_78 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_77;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_79 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_78;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_80 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_79;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_81 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_80;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_82 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_81;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_83 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_82;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_84 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_83;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_85 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_84;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_86 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_85;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_87 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_86;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_88 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_87;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_89 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_88;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_90 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_89;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_91 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_90;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_92 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_91;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_93 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_92;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_94 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_93;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_95 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_94;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_96 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_95;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_97 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_96;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_98 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_97;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_99 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_98;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_100 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_99;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_101 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_100;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_102 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_101;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_103 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_102;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_104 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_103;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_105 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_104;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_106 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_105;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_107 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_106;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_108 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_107;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_109 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_108;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_110 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_109;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_111 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_110;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_112 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_111;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_113 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_112;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_114 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_113;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_115 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_114;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_116 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_115;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_117 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_116;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_118 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_117;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_119 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_118;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_120 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_119;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_121 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_120;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_122 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_121;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_123 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_122;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_124 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_123;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_125 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_124;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_126 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_125;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_127 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_126;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_128 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_127;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_129 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_128;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_130 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_129;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_131 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_130;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_132 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_131;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_133 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_132;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_134 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_133;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_135 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_134;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_136 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_135;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_137 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_136;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_138 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_137;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_139 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_138;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_140 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_139;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_141 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_140;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_142 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_141;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_143 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_142;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_144 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_143;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_145 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_144;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_146 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_145;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_147 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_146;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_148 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_147;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_149 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_148;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_150 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_149;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_151 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_150;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_152 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_151;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_153 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_152;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_154 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_153;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_155 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_154;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_156 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_155;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_157 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_156;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_158 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_157;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_159 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_158;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_160 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_159;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_161 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_160;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_162 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_161;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_163 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_162;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_164 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_163;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_165 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_164;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_166 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_165;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_167 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_166;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_168 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_167;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_169 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_168;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_170 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_169;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_171 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_170;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_172 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_171;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_173 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_172;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_174 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_173;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_175 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_174;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_176 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_175;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_177 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_176;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_178 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_177;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_179 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_178;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_180 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_179;
      dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_181 <= dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51_stage_180;
      dark_weights_normed_gauss_blur_1_update_0_stage_77 <= dark_weights_normed_gauss_blur_1_update_0;
      dark_weights_normed_gauss_blur_1_update_0_stage_78 <= dark_weights_normed_gauss_blur_1_update_0_stage_77;
      dark_weights_normed_gauss_blur_1_update_0_stage_79 <= dark_weights_normed_gauss_blur_1_update_0_stage_78;
      dark_weights_normed_gauss_blur_1_update_0_stage_80 <= dark_weights_normed_gauss_blur_1_update_0_stage_79;
      dark_weights_normed_gauss_blur_1_update_0_stage_81 <= dark_weights_normed_gauss_blur_1_update_0_stage_80;
      dark_weights_normed_gauss_blur_1_update_0_stage_82 <= dark_weights_normed_gauss_blur_1_update_0_stage_81;
      dark_weights_normed_gauss_blur_1_update_0_stage_83 <= dark_weights_normed_gauss_blur_1_update_0_stage_82;
      dark_weights_normed_gauss_blur_1_update_0_stage_84 <= dark_weights_normed_gauss_blur_1_update_0_stage_83;
      dark_weights_normed_gauss_blur_1_update_0_stage_85 <= dark_weights_normed_gauss_blur_1_update_0_stage_84;
      dark_weights_normed_gauss_blur_1_update_0_stage_86 <= dark_weights_normed_gauss_blur_1_update_0_stage_85;
      dark_weights_normed_gauss_blur_1_update_0_stage_87 <= dark_weights_normed_gauss_blur_1_update_0_stage_86;
      dark_weights_normed_gauss_blur_1_update_0_stage_88 <= dark_weights_normed_gauss_blur_1_update_0_stage_87;
      dark_weights_normed_gauss_blur_1_update_0_stage_89 <= dark_weights_normed_gauss_blur_1_update_0_stage_88;
      dark_weights_normed_gauss_blur_1_update_0_stage_90 <= dark_weights_normed_gauss_blur_1_update_0_stage_89;
      dark_weights_normed_gauss_blur_1_update_0_stage_91 <= dark_weights_normed_gauss_blur_1_update_0_stage_90;
      dark_weights_normed_gauss_blur_1_update_0_stage_92 <= dark_weights_normed_gauss_blur_1_update_0_stage_91;
      dark_weights_normed_gauss_blur_1_update_0_stage_93 <= dark_weights_normed_gauss_blur_1_update_0_stage_92;
      dark_weights_normed_gauss_blur_1_update_0_stage_94 <= dark_weights_normed_gauss_blur_1_update_0_stage_93;
      dark_weights_normed_gauss_blur_1_update_0_stage_95 <= dark_weights_normed_gauss_blur_1_update_0_stage_94;
      dark_weights_normed_gauss_blur_1_update_0_stage_96 <= dark_weights_normed_gauss_blur_1_update_0_stage_95;
      dark_weights_normed_gauss_blur_1_update_0_stage_97 <= dark_weights_normed_gauss_blur_1_update_0_stage_96;
      dark_weights_normed_gauss_blur_1_update_0_stage_98 <= dark_weights_normed_gauss_blur_1_update_0_stage_97;
      dark_weights_normed_gauss_blur_1_update_0_stage_99 <= dark_weights_normed_gauss_blur_1_update_0_stage_98;
      dark_weights_normed_gauss_blur_1_update_0_stage_100 <= dark_weights_normed_gauss_blur_1_update_0_stage_99;
      dark_weights_normed_gauss_blur_1_update_0_stage_101 <= dark_weights_normed_gauss_blur_1_update_0_stage_100;
      dark_weights_normed_gauss_blur_1_update_0_stage_102 <= dark_weights_normed_gauss_blur_1_update_0_stage_101;
      dark_weights_normed_gauss_blur_1_update_0_stage_103 <= dark_weights_normed_gauss_blur_1_update_0_stage_102;
      dark_weights_normed_gauss_blur_1_update_0_stage_104 <= dark_weights_normed_gauss_blur_1_update_0_stage_103;
      dark_weights_normed_gauss_blur_1_update_0_stage_105 <= dark_weights_normed_gauss_blur_1_update_0_stage_104;
      dark_weights_normed_gauss_blur_1_update_0_stage_106 <= dark_weights_normed_gauss_blur_1_update_0_stage_105;
      dark_weights_normed_gauss_blur_1_update_0_stage_107 <= dark_weights_normed_gauss_blur_1_update_0_stage_106;
      dark_weights_normed_gauss_blur_1_update_0_stage_108 <= dark_weights_normed_gauss_blur_1_update_0_stage_107;
      dark_weights_normed_gauss_blur_1_update_0_stage_109 <= dark_weights_normed_gauss_blur_1_update_0_stage_108;
      dark_weights_normed_gauss_blur_1_update_0_stage_110 <= dark_weights_normed_gauss_blur_1_update_0_stage_109;
      dark_weights_normed_gauss_blur_1_update_0_stage_111 <= dark_weights_normed_gauss_blur_1_update_0_stage_110;
      dark_weights_normed_gauss_blur_1_update_0_stage_112 <= dark_weights_normed_gauss_blur_1_update_0_stage_111;
      dark_weights_normed_gauss_blur_1_update_0_stage_113 <= dark_weights_normed_gauss_blur_1_update_0_stage_112;
      dark_weights_normed_gauss_blur_1_update_0_stage_114 <= dark_weights_normed_gauss_blur_1_update_0_stage_113;
      dark_weights_normed_gauss_blur_1_update_0_stage_115 <= dark_weights_normed_gauss_blur_1_update_0_stage_114;
      dark_weights_normed_gauss_blur_1_update_0_stage_116 <= dark_weights_normed_gauss_blur_1_update_0_stage_115;
      dark_weights_normed_gauss_blur_1_update_0_stage_117 <= dark_weights_normed_gauss_blur_1_update_0_stage_116;
      dark_weights_normed_gauss_blur_1_update_0_stage_118 <= dark_weights_normed_gauss_blur_1_update_0_stage_117;
      dark_weights_normed_gauss_blur_1_update_0_stage_119 <= dark_weights_normed_gauss_blur_1_update_0_stage_118;
      dark_weights_normed_gauss_blur_1_update_0_stage_120 <= dark_weights_normed_gauss_blur_1_update_0_stage_119;
      dark_weights_normed_gauss_blur_1_update_0_stage_121 <= dark_weights_normed_gauss_blur_1_update_0_stage_120;
      dark_weights_normed_gauss_blur_1_update_0_stage_122 <= dark_weights_normed_gauss_blur_1_update_0_stage_121;
      dark_weights_normed_gauss_blur_1_update_0_stage_123 <= dark_weights_normed_gauss_blur_1_update_0_stage_122;
      dark_weights_normed_gauss_blur_1_update_0_stage_124 <= dark_weights_normed_gauss_blur_1_update_0_stage_123;
      dark_weights_normed_gauss_blur_1_update_0_stage_125 <= dark_weights_normed_gauss_blur_1_update_0_stage_124;
      dark_weights_normed_gauss_blur_1_update_0_stage_126 <= dark_weights_normed_gauss_blur_1_update_0_stage_125;
      dark_weights_normed_gauss_blur_1_update_0_stage_127 <= dark_weights_normed_gauss_blur_1_update_0_stage_126;
      dark_weights_normed_gauss_blur_1_update_0_stage_128 <= dark_weights_normed_gauss_blur_1_update_0_stage_127;
      dark_weights_normed_gauss_blur_1_update_0_stage_129 <= dark_weights_normed_gauss_blur_1_update_0_stage_128;
      dark_weights_normed_gauss_blur_1_update_0_stage_130 <= dark_weights_normed_gauss_blur_1_update_0_stage_129;
      dark_weights_normed_gauss_blur_1_update_0_stage_131 <= dark_weights_normed_gauss_blur_1_update_0_stage_130;
      dark_weights_normed_gauss_blur_1_update_0_stage_132 <= dark_weights_normed_gauss_blur_1_update_0_stage_131;
      dark_weights_normed_gauss_blur_1_update_0_stage_133 <= dark_weights_normed_gauss_blur_1_update_0_stage_132;
      dark_weights_normed_gauss_blur_1_update_0_stage_134 <= dark_weights_normed_gauss_blur_1_update_0_stage_133;
      dark_weights_normed_gauss_blur_1_update_0_stage_135 <= dark_weights_normed_gauss_blur_1_update_0_stage_134;
      dark_weights_normed_gauss_blur_1_update_0_stage_136 <= dark_weights_normed_gauss_blur_1_update_0_stage_135;
      dark_weights_normed_gauss_blur_1_update_0_stage_137 <= dark_weights_normed_gauss_blur_1_update_0_stage_136;
      dark_weights_normed_gauss_blur_1_update_0_stage_138 <= dark_weights_normed_gauss_blur_1_update_0_stage_137;
      dark_weights_normed_gauss_blur_1_update_0_stage_139 <= dark_weights_normed_gauss_blur_1_update_0_stage_138;
      dark_weights_normed_gauss_blur_1_update_0_stage_140 <= dark_weights_normed_gauss_blur_1_update_0_stage_139;
      dark_weights_normed_gauss_blur_1_update_0_stage_141 <= dark_weights_normed_gauss_blur_1_update_0_stage_140;
      dark_weights_normed_gauss_blur_1_update_0_stage_142 <= dark_weights_normed_gauss_blur_1_update_0_stage_141;
      dark_weights_normed_gauss_blur_1_update_0_stage_143 <= dark_weights_normed_gauss_blur_1_update_0_stage_142;
      dark_weights_normed_gauss_blur_1_update_0_stage_144 <= dark_weights_normed_gauss_blur_1_update_0_stage_143;
      dark_weights_normed_gauss_blur_1_update_0_stage_145 <= dark_weights_normed_gauss_blur_1_update_0_stage_144;
      dark_weights_normed_gauss_blur_1_update_0_stage_146 <= dark_weights_normed_gauss_blur_1_update_0_stage_145;
      dark_weights_normed_gauss_blur_1_update_0_stage_147 <= dark_weights_normed_gauss_blur_1_update_0_stage_146;
      dark_weights_normed_gauss_blur_1_update_0_stage_148 <= dark_weights_normed_gauss_blur_1_update_0_stage_147;
      dark_weights_normed_gauss_blur_1_update_0_stage_149 <= dark_weights_normed_gauss_blur_1_update_0_stage_148;
      dark_weights_normed_gauss_blur_1_update_0_stage_150 <= dark_weights_normed_gauss_blur_1_update_0_stage_149;
      dark_weights_normed_gauss_blur_1_update_0_stage_151 <= dark_weights_normed_gauss_blur_1_update_0_stage_150;
      dark_weights_normed_gauss_blur_1_update_0_stage_152 <= dark_weights_normed_gauss_blur_1_update_0_stage_151;
      dark_weights_normed_gauss_blur_1_update_0_stage_153 <= dark_weights_normed_gauss_blur_1_update_0_stage_152;
      dark_weights_normed_gauss_blur_1_update_0_stage_154 <= dark_weights_normed_gauss_blur_1_update_0_stage_153;
      dark_weights_normed_gauss_blur_1_update_0_stage_155 <= dark_weights_normed_gauss_blur_1_update_0_stage_154;
      dark_weights_normed_gauss_blur_1_update_0_stage_156 <= dark_weights_normed_gauss_blur_1_update_0_stage_155;
      dark_weights_normed_gauss_blur_1_update_0_stage_157 <= dark_weights_normed_gauss_blur_1_update_0_stage_156;
      dark_weights_normed_gauss_blur_1_update_0_stage_158 <= dark_weights_normed_gauss_blur_1_update_0_stage_157;
      dark_weights_normed_gauss_blur_1_update_0_stage_159 <= dark_weights_normed_gauss_blur_1_update_0_stage_158;
      dark_weights_normed_gauss_blur_1_update_0_stage_160 <= dark_weights_normed_gauss_blur_1_update_0_stage_159;
      dark_weights_normed_gauss_blur_1_update_0_stage_161 <= dark_weights_normed_gauss_blur_1_update_0_stage_160;
      dark_weights_normed_gauss_blur_1_update_0_stage_162 <= dark_weights_normed_gauss_blur_1_update_0_stage_161;
      dark_weights_normed_gauss_blur_1_update_0_stage_163 <= dark_weights_normed_gauss_blur_1_update_0_stage_162;
      dark_weights_normed_gauss_blur_1_update_0_stage_164 <= dark_weights_normed_gauss_blur_1_update_0_stage_163;
      dark_weights_normed_gauss_blur_1_update_0_stage_165 <= dark_weights_normed_gauss_blur_1_update_0_stage_164;
      dark_weights_normed_gauss_blur_1_update_0_stage_166 <= dark_weights_normed_gauss_blur_1_update_0_stage_165;
      dark_weights_normed_gauss_blur_1_update_0_stage_167 <= dark_weights_normed_gauss_blur_1_update_0_stage_166;
      dark_weights_normed_gauss_blur_1_update_0_stage_168 <= dark_weights_normed_gauss_blur_1_update_0_stage_167;
      dark_weights_normed_gauss_blur_1_update_0_stage_169 <= dark_weights_normed_gauss_blur_1_update_0_stage_168;
      dark_weights_normed_gauss_blur_1_update_0_stage_170 <= dark_weights_normed_gauss_blur_1_update_0_stage_169;
      dark_weights_normed_gauss_blur_1_update_0_stage_171 <= dark_weights_normed_gauss_blur_1_update_0_stage_170;
      dark_weights_normed_gauss_blur_1_update_0_stage_172 <= dark_weights_normed_gauss_blur_1_update_0_stage_171;
      dark_weights_normed_gauss_blur_1_update_0_stage_173 <= dark_weights_normed_gauss_blur_1_update_0_stage_172;
      dark_weights_normed_gauss_blur_1_update_0_stage_174 <= dark_weights_normed_gauss_blur_1_update_0_stage_173;
      dark_weights_normed_gauss_blur_1_update_0_stage_175 <= dark_weights_normed_gauss_blur_1_update_0_stage_174;
      dark_weights_normed_gauss_blur_1_update_0_stage_176 <= dark_weights_normed_gauss_blur_1_update_0_stage_175;
      dark_weights_normed_gauss_blur_1_update_0_stage_177 <= dark_weights_normed_gauss_blur_1_update_0_stage_176;
      dark_weights_normed_gauss_blur_1_update_0_stage_178 <= dark_weights_normed_gauss_blur_1_update_0_stage_177;
      dark_weights_normed_gauss_blur_1_update_0_stage_179 <= dark_weights_normed_gauss_blur_1_update_0_stage_178;
      dark_weights_normed_gauss_blur_1_update_0_stage_180 <= dark_weights_normed_gauss_blur_1_update_0_stage_179;
      dark_weights_normed_gauss_blur_1_update_0_stage_181 <= dark_weights_normed_gauss_blur_1_update_0_stage_180;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_78 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_79 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_78;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_80 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_79;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_81 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_80;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_82 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_81;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_83 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_82;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_84 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_83;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_85 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_84;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_86 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_85;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_87 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_86;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_88 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_87;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_89 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_88;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_90 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_89;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_91 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_90;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_92 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_91;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_93 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_92;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_94 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_93;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_95 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_94;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_96 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_95;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_97 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_96;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_98 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_97;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_99 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_98;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_100 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_99;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_101 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_100;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_102 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_101;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_103 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_102;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_104 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_103;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_105 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_104;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_106 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_105;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_107 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_106;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_108 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_107;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_109 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_108;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_110 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_109;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_111 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_110;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_112 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_111;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_113 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_112;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_114 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_113;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_115 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_114;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_116 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_115;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_117 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_116;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_118 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_117;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_119 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_118;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_120 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_119;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_121 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_120;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_122 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_121;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_123 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_122;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_124 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_123;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_125 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_124;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_126 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_125;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_127 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_126;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_128 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_127;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_129 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_128;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_130 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_129;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_131 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_130;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_132 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_131;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_133 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_132;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_134 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_133;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_135 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_134;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_136 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_135;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_137 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_136;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_138 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_137;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_139 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_138;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_140 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_139;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_141 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_140;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_142 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_141;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_143 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_142;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_144 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_143;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_145 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_144;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_146 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_145;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_147 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_146;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_148 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_147;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_149 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_148;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_150 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_149;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_151 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_150;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_152 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_151;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_153 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_152;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_154 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_153;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_155 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_154;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_156 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_155;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_157 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_156;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_158 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_157;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_159 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_158;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_160 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_159;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_161 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_160;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_162 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_161;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_163 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_162;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_164 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_163;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_165 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_164;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_166 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_165;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_167 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_166;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_168 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_167;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_169 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_168;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_170 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_169;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_171 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_170;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_172 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_171;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_173 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_172;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_174 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_173;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_175 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_174;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_176 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_175;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_177 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_176;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_178 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_177;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_179 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_178;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_180 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_179;
      dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_181 <= dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52_stage_180;
      dark_laplace_us_1_update_0_stage_92 <= dark_laplace_us_1_update_0;
      dark_laplace_us_1_update_0_stage_93 <= dark_laplace_us_1_update_0_stage_92;
      dark_laplace_us_1_update_0_stage_94 <= dark_laplace_us_1_update_0_stage_93;
      dark_laplace_us_1_update_0_stage_95 <= dark_laplace_us_1_update_0_stage_94;
      dark_laplace_us_1_update_0_stage_96 <= dark_laplace_us_1_update_0_stage_95;
      dark_laplace_us_1_update_0_stage_97 <= dark_laplace_us_1_update_0_stage_96;
      dark_laplace_us_1_update_0_stage_98 <= dark_laplace_us_1_update_0_stage_97;
      dark_laplace_us_1_update_0_stage_99 <= dark_laplace_us_1_update_0_stage_98;
      dark_laplace_us_1_update_0_stage_100 <= dark_laplace_us_1_update_0_stage_99;
      dark_laplace_us_1_update_0_stage_101 <= dark_laplace_us_1_update_0_stage_100;
      dark_laplace_us_1_update_0_stage_102 <= dark_laplace_us_1_update_0_stage_101;
      dark_laplace_us_1_update_0_stage_103 <= dark_laplace_us_1_update_0_stage_102;
      dark_laplace_us_1_update_0_stage_104 <= dark_laplace_us_1_update_0_stage_103;
      dark_laplace_us_1_update_0_stage_105 <= dark_laplace_us_1_update_0_stage_104;
      dark_laplace_us_1_update_0_stage_106 <= dark_laplace_us_1_update_0_stage_105;
      dark_laplace_us_1_update_0_stage_107 <= dark_laplace_us_1_update_0_stage_106;
      dark_laplace_us_1_update_0_stage_108 <= dark_laplace_us_1_update_0_stage_107;
      dark_laplace_us_1_update_0_stage_109 <= dark_laplace_us_1_update_0_stage_108;
      dark_laplace_us_1_update_0_stage_110 <= dark_laplace_us_1_update_0_stage_109;
      dark_laplace_us_1_update_0_stage_111 <= dark_laplace_us_1_update_0_stage_110;
      dark_laplace_us_1_update_0_stage_112 <= dark_laplace_us_1_update_0_stage_111;
      dark_laplace_us_1_update_0_stage_113 <= dark_laplace_us_1_update_0_stage_112;
      dark_laplace_us_1_update_0_stage_114 <= dark_laplace_us_1_update_0_stage_113;
      dark_laplace_us_1_update_0_stage_115 <= dark_laplace_us_1_update_0_stage_114;
      dark_laplace_us_1_update_0_stage_116 <= dark_laplace_us_1_update_0_stage_115;
      dark_laplace_us_1_update_0_stage_117 <= dark_laplace_us_1_update_0_stage_116;
      dark_laplace_us_1_update_0_stage_118 <= dark_laplace_us_1_update_0_stage_117;
      dark_laplace_us_1_update_0_stage_119 <= dark_laplace_us_1_update_0_stage_118;
      dark_laplace_us_1_update_0_stage_120 <= dark_laplace_us_1_update_0_stage_119;
      dark_laplace_us_1_update_0_stage_121 <= dark_laplace_us_1_update_0_stage_120;
      dark_laplace_us_1_update_0_stage_122 <= dark_laplace_us_1_update_0_stage_121;
      dark_laplace_us_1_update_0_stage_123 <= dark_laplace_us_1_update_0_stage_122;
      dark_laplace_us_1_update_0_stage_124 <= dark_laplace_us_1_update_0_stage_123;
      dark_laplace_us_1_update_0_stage_125 <= dark_laplace_us_1_update_0_stage_124;
      dark_laplace_us_1_update_0_stage_126 <= dark_laplace_us_1_update_0_stage_125;
      dark_laplace_us_1_update_0_stage_127 <= dark_laplace_us_1_update_0_stage_126;
      dark_laplace_us_1_update_0_stage_128 <= dark_laplace_us_1_update_0_stage_127;
      dark_laplace_us_1_update_0_stage_129 <= dark_laplace_us_1_update_0_stage_128;
      dark_laplace_us_1_update_0_stage_130 <= dark_laplace_us_1_update_0_stage_129;
      dark_laplace_us_1_update_0_stage_131 <= dark_laplace_us_1_update_0_stage_130;
      dark_laplace_us_1_update_0_stage_132 <= dark_laplace_us_1_update_0_stage_131;
      dark_laplace_us_1_update_0_stage_133 <= dark_laplace_us_1_update_0_stage_132;
      dark_laplace_us_1_update_0_stage_134 <= dark_laplace_us_1_update_0_stage_133;
      dark_laplace_us_1_update_0_stage_135 <= dark_laplace_us_1_update_0_stage_134;
      dark_laplace_us_1_update_0_stage_136 <= dark_laplace_us_1_update_0_stage_135;
      dark_laplace_us_1_update_0_stage_137 <= dark_laplace_us_1_update_0_stage_136;
      dark_laplace_us_1_update_0_stage_138 <= dark_laplace_us_1_update_0_stage_137;
      dark_laplace_us_1_update_0_stage_139 <= dark_laplace_us_1_update_0_stage_138;
      dark_laplace_us_1_update_0_stage_140 <= dark_laplace_us_1_update_0_stage_139;
      dark_laplace_us_1_update_0_stage_141 <= dark_laplace_us_1_update_0_stage_140;
      dark_laplace_us_1_update_0_stage_142 <= dark_laplace_us_1_update_0_stage_141;
      dark_laplace_us_1_update_0_stage_143 <= dark_laplace_us_1_update_0_stage_142;
      dark_laplace_us_1_update_0_stage_144 <= dark_laplace_us_1_update_0_stage_143;
      dark_laplace_us_1_update_0_stage_145 <= dark_laplace_us_1_update_0_stage_144;
      dark_laplace_us_1_update_0_stage_146 <= dark_laplace_us_1_update_0_stage_145;
      dark_laplace_us_1_update_0_stage_147 <= dark_laplace_us_1_update_0_stage_146;
      dark_laplace_us_1_update_0_stage_148 <= dark_laplace_us_1_update_0_stage_147;
      dark_laplace_us_1_update_0_stage_149 <= dark_laplace_us_1_update_0_stage_148;
      dark_laplace_us_1_update_0_stage_150 <= dark_laplace_us_1_update_0_stage_149;
      dark_laplace_us_1_update_0_stage_151 <= dark_laplace_us_1_update_0_stage_150;
      dark_laplace_us_1_update_0_stage_152 <= dark_laplace_us_1_update_0_stage_151;
      dark_laplace_us_1_update_0_stage_153 <= dark_laplace_us_1_update_0_stage_152;
      dark_laplace_us_1_update_0_stage_154 <= dark_laplace_us_1_update_0_stage_153;
      dark_laplace_us_1_update_0_stage_155 <= dark_laplace_us_1_update_0_stage_154;
      dark_laplace_us_1_update_0_stage_156 <= dark_laplace_us_1_update_0_stage_155;
      dark_laplace_us_1_update_0_stage_157 <= dark_laplace_us_1_update_0_stage_156;
      dark_laplace_us_1_update_0_stage_158 <= dark_laplace_us_1_update_0_stage_157;
      dark_laplace_us_1_update_0_stage_159 <= dark_laplace_us_1_update_0_stage_158;
      dark_laplace_us_1_update_0_stage_160 <= dark_laplace_us_1_update_0_stage_159;
      dark_laplace_us_1_update_0_stage_161 <= dark_laplace_us_1_update_0_stage_160;
      dark_laplace_us_1_update_0_stage_162 <= dark_laplace_us_1_update_0_stage_161;
      dark_laplace_us_1_update_0_stage_163 <= dark_laplace_us_1_update_0_stage_162;
      dark_laplace_us_1_update_0_stage_164 <= dark_laplace_us_1_update_0_stage_163;
      dark_laplace_us_1_update_0_stage_165 <= dark_laplace_us_1_update_0_stage_164;
      dark_laplace_us_1_update_0_stage_166 <= dark_laplace_us_1_update_0_stage_165;
      dark_laplace_us_1_update_0_stage_167 <= dark_laplace_us_1_update_0_stage_166;
      dark_laplace_us_1_update_0_stage_168 <= dark_laplace_us_1_update_0_stage_167;
      dark_laplace_us_1_update_0_stage_169 <= dark_laplace_us_1_update_0_stage_168;
      dark_laplace_us_1_update_0_stage_170 <= dark_laplace_us_1_update_0_stage_169;
      dark_laplace_us_1_update_0_stage_171 <= dark_laplace_us_1_update_0_stage_170;
      dark_laplace_us_1_update_0_stage_172 <= dark_laplace_us_1_update_0_stage_171;
      dark_laplace_us_1_update_0_stage_173 <= dark_laplace_us_1_update_0_stage_172;
      dark_laplace_us_1_update_0_stage_174 <= dark_laplace_us_1_update_0_stage_173;
      dark_laplace_us_1_update_0_stage_175 <= dark_laplace_us_1_update_0_stage_174;
      dark_laplace_us_1_update_0_stage_176 <= dark_laplace_us_1_update_0_stage_175;
      dark_laplace_us_1_update_0_stage_177 <= dark_laplace_us_1_update_0_stage_176;
      dark_laplace_us_1_update_0_stage_178 <= dark_laplace_us_1_update_0_stage_177;
      dark_laplace_us_1_update_0_stage_179 <= dark_laplace_us_1_update_0_stage_178;
      dark_laplace_us_1_update_0_stage_180 <= dark_laplace_us_1_update_0_stage_179;
      dark_laplace_us_1_update_0_stage_181 <= dark_laplace_us_1_update_0_stage_180;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_93 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_94 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_93;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_95 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_94;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_96 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_95;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_97 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_96;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_98 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_97;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_99 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_98;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_100 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_99;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_101 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_100;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_102 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_101;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_103 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_102;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_104 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_103;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_105 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_104;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_106 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_105;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_107 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_106;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_108 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_107;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_109 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_108;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_110 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_109;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_111 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_110;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_112 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_111;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_113 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_112;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_114 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_113;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_115 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_114;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_116 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_115;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_117 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_116;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_118 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_117;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_119 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_118;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_120 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_119;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_121 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_120;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_122 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_121;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_123 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_122;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_124 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_123;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_125 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_124;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_126 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_125;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_127 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_126;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_128 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_127;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_129 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_128;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_130 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_129;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_131 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_130;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_132 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_131;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_133 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_132;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_134 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_133;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_135 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_134;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_136 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_135;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_137 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_136;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_138 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_137;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_139 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_138;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_140 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_139;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_141 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_140;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_142 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_141;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_143 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_142;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_144 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_143;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_145 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_144;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_146 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_145;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_147 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_146;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_148 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_147;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_149 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_148;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_150 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_149;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_151 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_150;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_152 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_151;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_153 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_152;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_154 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_153;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_155 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_154;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_156 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_155;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_157 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_156;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_158 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_157;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_159 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_158;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_160 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_159;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_161 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_160;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_162 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_161;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_163 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_162;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_164 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_163;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_165 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_164;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_166 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_165;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_167 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_166;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_168 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_167;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_169 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_168;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_170 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_169;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_171 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_170;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_172 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_171;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_173 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_172;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_174 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_173;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_175 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_174;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_176 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_175;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_177 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_176;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_178 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_177;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_179 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_178;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_180 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_179;
      dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_181 <= dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62_stage_180;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_100 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_101 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_100;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_102 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_101;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_103 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_102;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_104 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_103;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_105 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_104;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_106 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_105;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_107 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_106;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_108 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_107;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_109 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_108;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_110 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_109;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_111 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_110;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_112 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_111;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_113 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_112;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_114 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_113;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_115 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_114;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_116 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_115;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_117 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_116;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_118 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_117;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_119 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_118;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_120 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_119;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_121 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_120;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_122 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_121;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_123 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_122;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_124 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_123;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_125 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_124;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_126 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_125;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_127 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_126;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_128 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_127;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_129 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_128;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_130 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_129;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_131 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_130;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_132 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_131;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_133 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_132;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_134 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_133;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_135 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_134;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_136 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_135;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_137 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_136;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_138 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_137;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_139 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_138;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_140 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_139;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_141 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_140;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_142 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_141;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_143 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_142;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_144 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_143;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_145 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_144;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_146 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_145;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_147 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_146;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_148 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_147;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_149 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_148;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_150 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_149;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_151 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_150;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_152 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_151;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_153 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_152;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_154 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_153;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_155 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_154;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_156 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_155;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_157 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_156;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_158 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_157;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_159 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_158;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_160 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_159;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_161 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_160;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_162 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_161;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_163 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_162;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_164 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_163;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_165 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_164;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_166 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_165;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_167 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_166;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_168 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_167;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_169 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_168;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_170 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_169;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_171 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_170;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_172 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_171;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_173 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_172;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_174 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_173;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_175 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_174;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_176 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_175;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_177 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_176;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_178 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_177;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_179 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_178;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_180 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_179;
      bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_181 <= bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67_stage_180;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_94 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_95 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_94;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_96 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_95;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_97 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_96;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_98 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_97;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_99 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_98;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_100 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_99;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_101 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_100;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_102 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_101;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_103 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_102;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_104 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_103;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_105 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_104;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_106 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_105;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_107 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_106;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_108 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_107;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_109 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_108;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_110 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_109;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_111 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_110;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_112 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_111;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_113 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_112;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_114 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_113;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_115 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_114;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_116 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_115;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_117 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_116;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_118 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_117;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_119 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_118;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_120 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_119;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_121 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_120;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_122 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_121;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_123 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_122;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_124 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_123;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_125 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_124;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_126 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_125;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_127 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_126;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_128 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_127;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_129 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_128;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_130 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_129;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_131 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_130;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_132 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_131;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_133 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_132;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_134 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_133;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_135 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_134;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_136 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_135;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_137 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_136;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_138 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_137;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_139 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_138;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_140 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_139;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_141 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_140;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_142 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_141;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_143 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_142;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_144 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_143;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_145 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_144;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_146 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_145;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_147 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_146;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_148 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_147;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_149 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_148;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_150 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_149;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_151 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_150;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_152 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_151;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_153 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_152;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_154 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_153;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_155 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_154;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_156 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_155;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_157 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_156;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_158 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_157;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_159 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_158;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_160 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_159;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_161 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_160;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_162 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_161;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_163 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_162;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_164 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_163;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_165 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_164;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_166 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_165;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_167 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_166;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_168 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_167;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_169 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_168;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_170 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_169;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_171 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_170;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_172 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_171;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_173 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_172;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_174 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_173;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_175 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_174;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_176 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_175;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_177 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_176;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_178 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_177;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_179 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_178;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_180 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_179;
      dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_181 <= dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63_stage_180;
      dark_weights_normed_gauss_ds_2_update_0_stage_95 <= dark_weights_normed_gauss_ds_2_update_0;
      dark_weights_normed_gauss_ds_2_update_0_stage_96 <= dark_weights_normed_gauss_ds_2_update_0_stage_95;
      dark_weights_normed_gauss_ds_2_update_0_stage_97 <= dark_weights_normed_gauss_ds_2_update_0_stage_96;
      dark_weights_normed_gauss_ds_2_update_0_stage_98 <= dark_weights_normed_gauss_ds_2_update_0_stage_97;
      dark_weights_normed_gauss_ds_2_update_0_stage_99 <= dark_weights_normed_gauss_ds_2_update_0_stage_98;
      dark_weights_normed_gauss_ds_2_update_0_stage_100 <= dark_weights_normed_gauss_ds_2_update_0_stage_99;
      dark_weights_normed_gauss_ds_2_update_0_stage_101 <= dark_weights_normed_gauss_ds_2_update_0_stage_100;
      dark_weights_normed_gauss_ds_2_update_0_stage_102 <= dark_weights_normed_gauss_ds_2_update_0_stage_101;
      dark_weights_normed_gauss_ds_2_update_0_stage_103 <= dark_weights_normed_gauss_ds_2_update_0_stage_102;
      dark_weights_normed_gauss_ds_2_update_0_stage_104 <= dark_weights_normed_gauss_ds_2_update_0_stage_103;
      dark_weights_normed_gauss_ds_2_update_0_stage_105 <= dark_weights_normed_gauss_ds_2_update_0_stage_104;
      dark_weights_normed_gauss_ds_2_update_0_stage_106 <= dark_weights_normed_gauss_ds_2_update_0_stage_105;
      dark_weights_normed_gauss_ds_2_update_0_stage_107 <= dark_weights_normed_gauss_ds_2_update_0_stage_106;
      dark_weights_normed_gauss_ds_2_update_0_stage_108 <= dark_weights_normed_gauss_ds_2_update_0_stage_107;
      dark_weights_normed_gauss_ds_2_update_0_stage_109 <= dark_weights_normed_gauss_ds_2_update_0_stage_108;
      dark_weights_normed_gauss_ds_2_update_0_stage_110 <= dark_weights_normed_gauss_ds_2_update_0_stage_109;
      dark_weights_normed_gauss_ds_2_update_0_stage_111 <= dark_weights_normed_gauss_ds_2_update_0_stage_110;
      dark_weights_normed_gauss_ds_2_update_0_stage_112 <= dark_weights_normed_gauss_ds_2_update_0_stage_111;
      dark_weights_normed_gauss_ds_2_update_0_stage_113 <= dark_weights_normed_gauss_ds_2_update_0_stage_112;
      dark_weights_normed_gauss_ds_2_update_0_stage_114 <= dark_weights_normed_gauss_ds_2_update_0_stage_113;
      dark_weights_normed_gauss_ds_2_update_0_stage_115 <= dark_weights_normed_gauss_ds_2_update_0_stage_114;
      dark_weights_normed_gauss_ds_2_update_0_stage_116 <= dark_weights_normed_gauss_ds_2_update_0_stage_115;
      dark_weights_normed_gauss_ds_2_update_0_stage_117 <= dark_weights_normed_gauss_ds_2_update_0_stage_116;
      dark_weights_normed_gauss_ds_2_update_0_stage_118 <= dark_weights_normed_gauss_ds_2_update_0_stage_117;
      dark_weights_normed_gauss_ds_2_update_0_stage_119 <= dark_weights_normed_gauss_ds_2_update_0_stage_118;
      dark_weights_normed_gauss_ds_2_update_0_stage_120 <= dark_weights_normed_gauss_ds_2_update_0_stage_119;
      dark_weights_normed_gauss_ds_2_update_0_stage_121 <= dark_weights_normed_gauss_ds_2_update_0_stage_120;
      dark_weights_normed_gauss_ds_2_update_0_stage_122 <= dark_weights_normed_gauss_ds_2_update_0_stage_121;
      dark_weights_normed_gauss_ds_2_update_0_stage_123 <= dark_weights_normed_gauss_ds_2_update_0_stage_122;
      dark_weights_normed_gauss_ds_2_update_0_stage_124 <= dark_weights_normed_gauss_ds_2_update_0_stage_123;
      dark_weights_normed_gauss_ds_2_update_0_stage_125 <= dark_weights_normed_gauss_ds_2_update_0_stage_124;
      dark_weights_normed_gauss_ds_2_update_0_stage_126 <= dark_weights_normed_gauss_ds_2_update_0_stage_125;
      dark_weights_normed_gauss_ds_2_update_0_stage_127 <= dark_weights_normed_gauss_ds_2_update_0_stage_126;
      dark_weights_normed_gauss_ds_2_update_0_stage_128 <= dark_weights_normed_gauss_ds_2_update_0_stage_127;
      dark_weights_normed_gauss_ds_2_update_0_stage_129 <= dark_weights_normed_gauss_ds_2_update_0_stage_128;
      dark_weights_normed_gauss_ds_2_update_0_stage_130 <= dark_weights_normed_gauss_ds_2_update_0_stage_129;
      dark_weights_normed_gauss_ds_2_update_0_stage_131 <= dark_weights_normed_gauss_ds_2_update_0_stage_130;
      dark_weights_normed_gauss_ds_2_update_0_stage_132 <= dark_weights_normed_gauss_ds_2_update_0_stage_131;
      dark_weights_normed_gauss_ds_2_update_0_stage_133 <= dark_weights_normed_gauss_ds_2_update_0_stage_132;
      dark_weights_normed_gauss_ds_2_update_0_stage_134 <= dark_weights_normed_gauss_ds_2_update_0_stage_133;
      dark_weights_normed_gauss_ds_2_update_0_stage_135 <= dark_weights_normed_gauss_ds_2_update_0_stage_134;
      dark_weights_normed_gauss_ds_2_update_0_stage_136 <= dark_weights_normed_gauss_ds_2_update_0_stage_135;
      dark_weights_normed_gauss_ds_2_update_0_stage_137 <= dark_weights_normed_gauss_ds_2_update_0_stage_136;
      dark_weights_normed_gauss_ds_2_update_0_stage_138 <= dark_weights_normed_gauss_ds_2_update_0_stage_137;
      dark_weights_normed_gauss_ds_2_update_0_stage_139 <= dark_weights_normed_gauss_ds_2_update_0_stage_138;
      dark_weights_normed_gauss_ds_2_update_0_stage_140 <= dark_weights_normed_gauss_ds_2_update_0_stage_139;
      dark_weights_normed_gauss_ds_2_update_0_stage_141 <= dark_weights_normed_gauss_ds_2_update_0_stage_140;
      dark_weights_normed_gauss_ds_2_update_0_stage_142 <= dark_weights_normed_gauss_ds_2_update_0_stage_141;
      dark_weights_normed_gauss_ds_2_update_0_stage_143 <= dark_weights_normed_gauss_ds_2_update_0_stage_142;
      dark_weights_normed_gauss_ds_2_update_0_stage_144 <= dark_weights_normed_gauss_ds_2_update_0_stage_143;
      dark_weights_normed_gauss_ds_2_update_0_stage_145 <= dark_weights_normed_gauss_ds_2_update_0_stage_144;
      dark_weights_normed_gauss_ds_2_update_0_stage_146 <= dark_weights_normed_gauss_ds_2_update_0_stage_145;
      dark_weights_normed_gauss_ds_2_update_0_stage_147 <= dark_weights_normed_gauss_ds_2_update_0_stage_146;
      dark_weights_normed_gauss_ds_2_update_0_stage_148 <= dark_weights_normed_gauss_ds_2_update_0_stage_147;
      dark_weights_normed_gauss_ds_2_update_0_stage_149 <= dark_weights_normed_gauss_ds_2_update_0_stage_148;
      dark_weights_normed_gauss_ds_2_update_0_stage_150 <= dark_weights_normed_gauss_ds_2_update_0_stage_149;
      dark_weights_normed_gauss_ds_2_update_0_stage_151 <= dark_weights_normed_gauss_ds_2_update_0_stage_150;
      dark_weights_normed_gauss_ds_2_update_0_stage_152 <= dark_weights_normed_gauss_ds_2_update_0_stage_151;
      dark_weights_normed_gauss_ds_2_update_0_stage_153 <= dark_weights_normed_gauss_ds_2_update_0_stage_152;
      dark_weights_normed_gauss_ds_2_update_0_stage_154 <= dark_weights_normed_gauss_ds_2_update_0_stage_153;
      dark_weights_normed_gauss_ds_2_update_0_stage_155 <= dark_weights_normed_gauss_ds_2_update_0_stage_154;
      dark_weights_normed_gauss_ds_2_update_0_stage_156 <= dark_weights_normed_gauss_ds_2_update_0_stage_155;
      dark_weights_normed_gauss_ds_2_update_0_stage_157 <= dark_weights_normed_gauss_ds_2_update_0_stage_156;
      dark_weights_normed_gauss_ds_2_update_0_stage_158 <= dark_weights_normed_gauss_ds_2_update_0_stage_157;
      dark_weights_normed_gauss_ds_2_update_0_stage_159 <= dark_weights_normed_gauss_ds_2_update_0_stage_158;
      dark_weights_normed_gauss_ds_2_update_0_stage_160 <= dark_weights_normed_gauss_ds_2_update_0_stage_159;
      dark_weights_normed_gauss_ds_2_update_0_stage_161 <= dark_weights_normed_gauss_ds_2_update_0_stage_160;
      dark_weights_normed_gauss_ds_2_update_0_stage_162 <= dark_weights_normed_gauss_ds_2_update_0_stage_161;
      dark_weights_normed_gauss_ds_2_update_0_stage_163 <= dark_weights_normed_gauss_ds_2_update_0_stage_162;
      dark_weights_normed_gauss_ds_2_update_0_stage_164 <= dark_weights_normed_gauss_ds_2_update_0_stage_163;
      dark_weights_normed_gauss_ds_2_update_0_stage_165 <= dark_weights_normed_gauss_ds_2_update_0_stage_164;
      dark_weights_normed_gauss_ds_2_update_0_stage_166 <= dark_weights_normed_gauss_ds_2_update_0_stage_165;
      dark_weights_normed_gauss_ds_2_update_0_stage_167 <= dark_weights_normed_gauss_ds_2_update_0_stage_166;
      dark_weights_normed_gauss_ds_2_update_0_stage_168 <= dark_weights_normed_gauss_ds_2_update_0_stage_167;
      dark_weights_normed_gauss_ds_2_update_0_stage_169 <= dark_weights_normed_gauss_ds_2_update_0_stage_168;
      dark_weights_normed_gauss_ds_2_update_0_stage_170 <= dark_weights_normed_gauss_ds_2_update_0_stage_169;
      dark_weights_normed_gauss_ds_2_update_0_stage_171 <= dark_weights_normed_gauss_ds_2_update_0_stage_170;
      dark_weights_normed_gauss_ds_2_update_0_stage_172 <= dark_weights_normed_gauss_ds_2_update_0_stage_171;
      dark_weights_normed_gauss_ds_2_update_0_stage_173 <= dark_weights_normed_gauss_ds_2_update_0_stage_172;
      dark_weights_normed_gauss_ds_2_update_0_stage_174 <= dark_weights_normed_gauss_ds_2_update_0_stage_173;
      dark_weights_normed_gauss_ds_2_update_0_stage_175 <= dark_weights_normed_gauss_ds_2_update_0_stage_174;
      dark_weights_normed_gauss_ds_2_update_0_stage_176 <= dark_weights_normed_gauss_ds_2_update_0_stage_175;
      dark_weights_normed_gauss_ds_2_update_0_stage_177 <= dark_weights_normed_gauss_ds_2_update_0_stage_176;
      dark_weights_normed_gauss_ds_2_update_0_stage_178 <= dark_weights_normed_gauss_ds_2_update_0_stage_177;
      dark_weights_normed_gauss_ds_2_update_0_stage_179 <= dark_weights_normed_gauss_ds_2_update_0_stage_178;
      dark_weights_normed_gauss_ds_2_update_0_stage_180 <= dark_weights_normed_gauss_ds_2_update_0_stage_179;
      dark_weights_normed_gauss_ds_2_update_0_stage_181 <= dark_weights_normed_gauss_ds_2_update_0_stage_180;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_96 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_97 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_96;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_98 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_97;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_99 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_98;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_100 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_99;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_101 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_100;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_102 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_101;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_103 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_102;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_104 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_103;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_105 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_104;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_106 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_105;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_107 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_106;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_108 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_107;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_109 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_108;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_110 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_109;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_111 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_110;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_112 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_111;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_113 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_112;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_114 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_113;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_115 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_114;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_116 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_115;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_117 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_116;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_118 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_117;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_119 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_118;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_120 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_119;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_121 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_120;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_122 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_121;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_123 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_122;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_124 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_123;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_125 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_124;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_126 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_125;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_127 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_126;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_128 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_127;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_129 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_128;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_130 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_129;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_131 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_130;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_132 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_131;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_133 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_132;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_134 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_133;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_135 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_134;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_136 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_135;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_137 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_136;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_138 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_137;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_139 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_138;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_140 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_139;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_141 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_140;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_142 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_141;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_143 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_142;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_144 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_143;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_145 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_144;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_146 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_145;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_147 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_146;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_148 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_147;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_149 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_148;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_150 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_149;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_151 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_150;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_152 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_151;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_153 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_152;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_154 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_153;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_155 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_154;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_156 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_155;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_157 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_156;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_158 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_157;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_159 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_158;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_160 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_159;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_161 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_160;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_162 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_161;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_163 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_162;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_164 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_163;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_165 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_164;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_166 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_165;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_167 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_166;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_168 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_167;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_169 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_168;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_170 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_169;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_171 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_170;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_172 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_171;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_173 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_172;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_174 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_173;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_175 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_174;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_176 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_175;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_177 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_176;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_178 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_177;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_179 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_178;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_180 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_179;
      dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_181 <= dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64_stage_180;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_101 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_102 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_101;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_103 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_102;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_104 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_103;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_105 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_104;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_106 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_105;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_107 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_106;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_108 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_107;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_109 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_108;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_110 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_109;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_111 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_110;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_112 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_111;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_113 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_112;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_114 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_113;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_115 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_114;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_116 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_115;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_117 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_116;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_118 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_117;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_119 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_118;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_120 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_119;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_121 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_120;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_122 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_121;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_123 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_122;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_124 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_123;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_125 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_124;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_126 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_125;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_127 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_126;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_128 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_127;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_129 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_128;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_130 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_129;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_131 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_130;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_132 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_131;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_133 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_132;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_134 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_133;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_135 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_134;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_136 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_135;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_137 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_136;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_138 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_137;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_139 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_138;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_140 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_139;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_141 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_140;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_142 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_141;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_143 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_142;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_144 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_143;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_145 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_144;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_146 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_145;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_147 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_146;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_148 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_147;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_149 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_148;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_150 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_149;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_151 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_150;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_152 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_151;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_153 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_152;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_154 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_153;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_155 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_154;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_156 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_155;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_157 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_156;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_158 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_157;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_159 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_158;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_160 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_159;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_161 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_160;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_162 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_161;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_163 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_162;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_164 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_163;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_165 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_164;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_166 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_165;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_167 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_166;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_168 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_167;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_169 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_168;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_170 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_169;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_171 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_170;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_172 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_171;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_173 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_172;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_174 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_173;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_175 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_174;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_176 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_175;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_177 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_176;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_178 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_177;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_179 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_178;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_180 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_179;
      bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_181 <= bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68_stage_180;
      bright_laplace_diff_1_update_0_stage_102 <= bright_laplace_diff_1_update_0;
      bright_laplace_diff_1_update_0_stage_103 <= bright_laplace_diff_1_update_0_stage_102;
      bright_laplace_diff_1_update_0_stage_104 <= bright_laplace_diff_1_update_0_stage_103;
      bright_laplace_diff_1_update_0_stage_105 <= bright_laplace_diff_1_update_0_stage_104;
      bright_laplace_diff_1_update_0_stage_106 <= bright_laplace_diff_1_update_0_stage_105;
      bright_laplace_diff_1_update_0_stage_107 <= bright_laplace_diff_1_update_0_stage_106;
      bright_laplace_diff_1_update_0_stage_108 <= bright_laplace_diff_1_update_0_stage_107;
      bright_laplace_diff_1_update_0_stage_109 <= bright_laplace_diff_1_update_0_stage_108;
      bright_laplace_diff_1_update_0_stage_110 <= bright_laplace_diff_1_update_0_stage_109;
      bright_laplace_diff_1_update_0_stage_111 <= bright_laplace_diff_1_update_0_stage_110;
      bright_laplace_diff_1_update_0_stage_112 <= bright_laplace_diff_1_update_0_stage_111;
      bright_laplace_diff_1_update_0_stage_113 <= bright_laplace_diff_1_update_0_stage_112;
      bright_laplace_diff_1_update_0_stage_114 <= bright_laplace_diff_1_update_0_stage_113;
      bright_laplace_diff_1_update_0_stage_115 <= bright_laplace_diff_1_update_0_stage_114;
      bright_laplace_diff_1_update_0_stage_116 <= bright_laplace_diff_1_update_0_stage_115;
      bright_laplace_diff_1_update_0_stage_117 <= bright_laplace_diff_1_update_0_stage_116;
      bright_laplace_diff_1_update_0_stage_118 <= bright_laplace_diff_1_update_0_stage_117;
      bright_laplace_diff_1_update_0_stage_119 <= bright_laplace_diff_1_update_0_stage_118;
      bright_laplace_diff_1_update_0_stage_120 <= bright_laplace_diff_1_update_0_stage_119;
      bright_laplace_diff_1_update_0_stage_121 <= bright_laplace_diff_1_update_0_stage_120;
      bright_laplace_diff_1_update_0_stage_122 <= bright_laplace_diff_1_update_0_stage_121;
      bright_laplace_diff_1_update_0_stage_123 <= bright_laplace_diff_1_update_0_stage_122;
      bright_laplace_diff_1_update_0_stage_124 <= bright_laplace_diff_1_update_0_stage_123;
      bright_laplace_diff_1_update_0_stage_125 <= bright_laplace_diff_1_update_0_stage_124;
      bright_laplace_diff_1_update_0_stage_126 <= bright_laplace_diff_1_update_0_stage_125;
      bright_laplace_diff_1_update_0_stage_127 <= bright_laplace_diff_1_update_0_stage_126;
      bright_laplace_diff_1_update_0_stage_128 <= bright_laplace_diff_1_update_0_stage_127;
      bright_laplace_diff_1_update_0_stage_129 <= bright_laplace_diff_1_update_0_stage_128;
      bright_laplace_diff_1_update_0_stage_130 <= bright_laplace_diff_1_update_0_stage_129;
      bright_laplace_diff_1_update_0_stage_131 <= bright_laplace_diff_1_update_0_stage_130;
      bright_laplace_diff_1_update_0_stage_132 <= bright_laplace_diff_1_update_0_stage_131;
      bright_laplace_diff_1_update_0_stage_133 <= bright_laplace_diff_1_update_0_stage_132;
      bright_laplace_diff_1_update_0_stage_134 <= bright_laplace_diff_1_update_0_stage_133;
      bright_laplace_diff_1_update_0_stage_135 <= bright_laplace_diff_1_update_0_stage_134;
      bright_laplace_diff_1_update_0_stage_136 <= bright_laplace_diff_1_update_0_stage_135;
      bright_laplace_diff_1_update_0_stage_137 <= bright_laplace_diff_1_update_0_stage_136;
      bright_laplace_diff_1_update_0_stage_138 <= bright_laplace_diff_1_update_0_stage_137;
      bright_laplace_diff_1_update_0_stage_139 <= bright_laplace_diff_1_update_0_stage_138;
      bright_laplace_diff_1_update_0_stage_140 <= bright_laplace_diff_1_update_0_stage_139;
      bright_laplace_diff_1_update_0_stage_141 <= bright_laplace_diff_1_update_0_stage_140;
      bright_laplace_diff_1_update_0_stage_142 <= bright_laplace_diff_1_update_0_stage_141;
      bright_laplace_diff_1_update_0_stage_143 <= bright_laplace_diff_1_update_0_stage_142;
      bright_laplace_diff_1_update_0_stage_144 <= bright_laplace_diff_1_update_0_stage_143;
      bright_laplace_diff_1_update_0_stage_145 <= bright_laplace_diff_1_update_0_stage_144;
      bright_laplace_diff_1_update_0_stage_146 <= bright_laplace_diff_1_update_0_stage_145;
      bright_laplace_diff_1_update_0_stage_147 <= bright_laplace_diff_1_update_0_stage_146;
      bright_laplace_diff_1_update_0_stage_148 <= bright_laplace_diff_1_update_0_stage_147;
      bright_laplace_diff_1_update_0_stage_149 <= bright_laplace_diff_1_update_0_stage_148;
      bright_laplace_diff_1_update_0_stage_150 <= bright_laplace_diff_1_update_0_stage_149;
      bright_laplace_diff_1_update_0_stage_151 <= bright_laplace_diff_1_update_0_stage_150;
      bright_laplace_diff_1_update_0_stage_152 <= bright_laplace_diff_1_update_0_stage_151;
      bright_laplace_diff_1_update_0_stage_153 <= bright_laplace_diff_1_update_0_stage_152;
      bright_laplace_diff_1_update_0_stage_154 <= bright_laplace_diff_1_update_0_stage_153;
      bright_laplace_diff_1_update_0_stage_155 <= bright_laplace_diff_1_update_0_stage_154;
      bright_laplace_diff_1_update_0_stage_156 <= bright_laplace_diff_1_update_0_stage_155;
      bright_laplace_diff_1_update_0_stage_157 <= bright_laplace_diff_1_update_0_stage_156;
      bright_laplace_diff_1_update_0_stage_158 <= bright_laplace_diff_1_update_0_stage_157;
      bright_laplace_diff_1_update_0_stage_159 <= bright_laplace_diff_1_update_0_stage_158;
      bright_laplace_diff_1_update_0_stage_160 <= bright_laplace_diff_1_update_0_stage_159;
      bright_laplace_diff_1_update_0_stage_161 <= bright_laplace_diff_1_update_0_stage_160;
      bright_laplace_diff_1_update_0_stage_162 <= bright_laplace_diff_1_update_0_stage_161;
      bright_laplace_diff_1_update_0_stage_163 <= bright_laplace_diff_1_update_0_stage_162;
      bright_laplace_diff_1_update_0_stage_164 <= bright_laplace_diff_1_update_0_stage_163;
      bright_laplace_diff_1_update_0_stage_165 <= bright_laplace_diff_1_update_0_stage_164;
      bright_laplace_diff_1_update_0_stage_166 <= bright_laplace_diff_1_update_0_stage_165;
      bright_laplace_diff_1_update_0_stage_167 <= bright_laplace_diff_1_update_0_stage_166;
      bright_laplace_diff_1_update_0_stage_168 <= bright_laplace_diff_1_update_0_stage_167;
      bright_laplace_diff_1_update_0_stage_169 <= bright_laplace_diff_1_update_0_stage_168;
      bright_laplace_diff_1_update_0_stage_170 <= bright_laplace_diff_1_update_0_stage_169;
      bright_laplace_diff_1_update_0_stage_171 <= bright_laplace_diff_1_update_0_stage_170;
      bright_laplace_diff_1_update_0_stage_172 <= bright_laplace_diff_1_update_0_stage_171;
      bright_laplace_diff_1_update_0_stage_173 <= bright_laplace_diff_1_update_0_stage_172;
      bright_laplace_diff_1_update_0_stage_174 <= bright_laplace_diff_1_update_0_stage_173;
      bright_laplace_diff_1_update_0_stage_175 <= bright_laplace_diff_1_update_0_stage_174;
      bright_laplace_diff_1_update_0_stage_176 <= bright_laplace_diff_1_update_0_stage_175;
      bright_laplace_diff_1_update_0_stage_177 <= bright_laplace_diff_1_update_0_stage_176;
      bright_laplace_diff_1_update_0_stage_178 <= bright_laplace_diff_1_update_0_stage_177;
      bright_laplace_diff_1_update_0_stage_179 <= bright_laplace_diff_1_update_0_stage_178;
      bright_laplace_diff_1_update_0_stage_180 <= bright_laplace_diff_1_update_0_stage_179;
      bright_laplace_diff_1_update_0_stage_181 <= bright_laplace_diff_1_update_0_stage_180;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_103 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_104 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_103;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_105 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_104;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_106 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_105;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_107 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_106;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_108 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_107;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_109 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_108;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_110 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_109;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_111 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_110;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_112 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_111;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_113 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_112;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_114 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_113;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_115 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_114;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_116 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_115;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_117 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_116;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_118 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_117;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_119 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_118;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_120 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_119;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_121 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_120;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_122 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_121;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_123 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_122;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_124 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_123;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_125 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_124;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_126 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_125;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_127 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_126;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_128 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_127;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_129 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_128;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_130 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_129;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_131 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_130;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_132 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_131;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_133 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_132;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_134 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_133;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_135 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_134;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_136 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_135;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_137 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_136;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_138 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_137;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_139 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_138;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_140 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_139;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_141 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_140;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_142 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_141;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_143 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_142;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_144 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_143;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_145 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_144;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_146 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_145;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_147 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_146;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_148 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_147;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_149 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_148;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_150 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_149;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_151 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_150;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_152 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_151;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_153 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_152;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_154 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_153;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_155 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_154;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_156 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_155;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_157 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_156;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_158 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_157;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_159 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_158;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_160 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_159;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_161 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_160;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_162 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_161;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_163 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_162;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_164 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_163;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_165 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_164;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_166 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_165;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_167 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_166;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_168 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_167;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_169 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_168;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_170 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_169;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_171 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_170;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_172 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_171;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_173 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_172;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_174 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_173;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_175 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_174;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_176 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_175;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_177 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_176;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_178 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_177;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_179 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_178;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_180 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_179;
      bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_181 <= bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69_stage_180;
      dark_weights_normed_gauss_blur_3_update_0_stage_108 <= dark_weights_normed_gauss_blur_3_update_0;
      dark_weights_normed_gauss_blur_3_update_0_stage_109 <= dark_weights_normed_gauss_blur_3_update_0_stage_108;
      dark_weights_normed_gauss_blur_3_update_0_stage_110 <= dark_weights_normed_gauss_blur_3_update_0_stage_109;
      dark_weights_normed_gauss_blur_3_update_0_stage_111 <= dark_weights_normed_gauss_blur_3_update_0_stage_110;
      dark_weights_normed_gauss_blur_3_update_0_stage_112 <= dark_weights_normed_gauss_blur_3_update_0_stage_111;
      dark_weights_normed_gauss_blur_3_update_0_stage_113 <= dark_weights_normed_gauss_blur_3_update_0_stage_112;
      dark_weights_normed_gauss_blur_3_update_0_stage_114 <= dark_weights_normed_gauss_blur_3_update_0_stage_113;
      dark_weights_normed_gauss_blur_3_update_0_stage_115 <= dark_weights_normed_gauss_blur_3_update_0_stage_114;
      dark_weights_normed_gauss_blur_3_update_0_stage_116 <= dark_weights_normed_gauss_blur_3_update_0_stage_115;
      dark_weights_normed_gauss_blur_3_update_0_stage_117 <= dark_weights_normed_gauss_blur_3_update_0_stage_116;
      dark_weights_normed_gauss_blur_3_update_0_stage_118 <= dark_weights_normed_gauss_blur_3_update_0_stage_117;
      dark_weights_normed_gauss_blur_3_update_0_stage_119 <= dark_weights_normed_gauss_blur_3_update_0_stage_118;
      dark_weights_normed_gauss_blur_3_update_0_stage_120 <= dark_weights_normed_gauss_blur_3_update_0_stage_119;
      dark_weights_normed_gauss_blur_3_update_0_stage_121 <= dark_weights_normed_gauss_blur_3_update_0_stage_120;
      dark_weights_normed_gauss_blur_3_update_0_stage_122 <= dark_weights_normed_gauss_blur_3_update_0_stage_121;
      dark_weights_normed_gauss_blur_3_update_0_stage_123 <= dark_weights_normed_gauss_blur_3_update_0_stage_122;
      dark_weights_normed_gauss_blur_3_update_0_stage_124 <= dark_weights_normed_gauss_blur_3_update_0_stage_123;
      dark_weights_normed_gauss_blur_3_update_0_stage_125 <= dark_weights_normed_gauss_blur_3_update_0_stage_124;
      dark_weights_normed_gauss_blur_3_update_0_stage_126 <= dark_weights_normed_gauss_blur_3_update_0_stage_125;
      dark_weights_normed_gauss_blur_3_update_0_stage_127 <= dark_weights_normed_gauss_blur_3_update_0_stage_126;
      dark_weights_normed_gauss_blur_3_update_0_stage_128 <= dark_weights_normed_gauss_blur_3_update_0_stage_127;
      dark_weights_normed_gauss_blur_3_update_0_stage_129 <= dark_weights_normed_gauss_blur_3_update_0_stage_128;
      dark_weights_normed_gauss_blur_3_update_0_stage_130 <= dark_weights_normed_gauss_blur_3_update_0_stage_129;
      dark_weights_normed_gauss_blur_3_update_0_stage_131 <= dark_weights_normed_gauss_blur_3_update_0_stage_130;
      dark_weights_normed_gauss_blur_3_update_0_stage_132 <= dark_weights_normed_gauss_blur_3_update_0_stage_131;
      dark_weights_normed_gauss_blur_3_update_0_stage_133 <= dark_weights_normed_gauss_blur_3_update_0_stage_132;
      dark_weights_normed_gauss_blur_3_update_0_stage_134 <= dark_weights_normed_gauss_blur_3_update_0_stage_133;
      dark_weights_normed_gauss_blur_3_update_0_stage_135 <= dark_weights_normed_gauss_blur_3_update_0_stage_134;
      dark_weights_normed_gauss_blur_3_update_0_stage_136 <= dark_weights_normed_gauss_blur_3_update_0_stage_135;
      dark_weights_normed_gauss_blur_3_update_0_stage_137 <= dark_weights_normed_gauss_blur_3_update_0_stage_136;
      dark_weights_normed_gauss_blur_3_update_0_stage_138 <= dark_weights_normed_gauss_blur_3_update_0_stage_137;
      dark_weights_normed_gauss_blur_3_update_0_stage_139 <= dark_weights_normed_gauss_blur_3_update_0_stage_138;
      dark_weights_normed_gauss_blur_3_update_0_stage_140 <= dark_weights_normed_gauss_blur_3_update_0_stage_139;
      dark_weights_normed_gauss_blur_3_update_0_stage_141 <= dark_weights_normed_gauss_blur_3_update_0_stage_140;
      dark_weights_normed_gauss_blur_3_update_0_stage_142 <= dark_weights_normed_gauss_blur_3_update_0_stage_141;
      dark_weights_normed_gauss_blur_3_update_0_stage_143 <= dark_weights_normed_gauss_blur_3_update_0_stage_142;
      dark_weights_normed_gauss_blur_3_update_0_stage_144 <= dark_weights_normed_gauss_blur_3_update_0_stage_143;
      dark_weights_normed_gauss_blur_3_update_0_stage_145 <= dark_weights_normed_gauss_blur_3_update_0_stage_144;
      dark_weights_normed_gauss_blur_3_update_0_stage_146 <= dark_weights_normed_gauss_blur_3_update_0_stage_145;
      dark_weights_normed_gauss_blur_3_update_0_stage_147 <= dark_weights_normed_gauss_blur_3_update_0_stage_146;
      dark_weights_normed_gauss_blur_3_update_0_stage_148 <= dark_weights_normed_gauss_blur_3_update_0_stage_147;
      dark_weights_normed_gauss_blur_3_update_0_stage_149 <= dark_weights_normed_gauss_blur_3_update_0_stage_148;
      dark_weights_normed_gauss_blur_3_update_0_stage_150 <= dark_weights_normed_gauss_blur_3_update_0_stage_149;
      dark_weights_normed_gauss_blur_3_update_0_stage_151 <= dark_weights_normed_gauss_blur_3_update_0_stage_150;
      dark_weights_normed_gauss_blur_3_update_0_stage_152 <= dark_weights_normed_gauss_blur_3_update_0_stage_151;
      dark_weights_normed_gauss_blur_3_update_0_stage_153 <= dark_weights_normed_gauss_blur_3_update_0_stage_152;
      dark_weights_normed_gauss_blur_3_update_0_stage_154 <= dark_weights_normed_gauss_blur_3_update_0_stage_153;
      dark_weights_normed_gauss_blur_3_update_0_stage_155 <= dark_weights_normed_gauss_blur_3_update_0_stage_154;
      dark_weights_normed_gauss_blur_3_update_0_stage_156 <= dark_weights_normed_gauss_blur_3_update_0_stage_155;
      dark_weights_normed_gauss_blur_3_update_0_stage_157 <= dark_weights_normed_gauss_blur_3_update_0_stage_156;
      dark_weights_normed_gauss_blur_3_update_0_stage_158 <= dark_weights_normed_gauss_blur_3_update_0_stage_157;
      dark_weights_normed_gauss_blur_3_update_0_stage_159 <= dark_weights_normed_gauss_blur_3_update_0_stage_158;
      dark_weights_normed_gauss_blur_3_update_0_stage_160 <= dark_weights_normed_gauss_blur_3_update_0_stage_159;
      dark_weights_normed_gauss_blur_3_update_0_stage_161 <= dark_weights_normed_gauss_blur_3_update_0_stage_160;
      dark_weights_normed_gauss_blur_3_update_0_stage_162 <= dark_weights_normed_gauss_blur_3_update_0_stage_161;
      dark_weights_normed_gauss_blur_3_update_0_stage_163 <= dark_weights_normed_gauss_blur_3_update_0_stage_162;
      dark_weights_normed_gauss_blur_3_update_0_stage_164 <= dark_weights_normed_gauss_blur_3_update_0_stage_163;
      dark_weights_normed_gauss_blur_3_update_0_stage_165 <= dark_weights_normed_gauss_blur_3_update_0_stage_164;
      dark_weights_normed_gauss_blur_3_update_0_stage_166 <= dark_weights_normed_gauss_blur_3_update_0_stage_165;
      dark_weights_normed_gauss_blur_3_update_0_stage_167 <= dark_weights_normed_gauss_blur_3_update_0_stage_166;
      dark_weights_normed_gauss_blur_3_update_0_stage_168 <= dark_weights_normed_gauss_blur_3_update_0_stage_167;
      dark_weights_normed_gauss_blur_3_update_0_stage_169 <= dark_weights_normed_gauss_blur_3_update_0_stage_168;
      dark_weights_normed_gauss_blur_3_update_0_stage_170 <= dark_weights_normed_gauss_blur_3_update_0_stage_169;
      dark_weights_normed_gauss_blur_3_update_0_stage_171 <= dark_weights_normed_gauss_blur_3_update_0_stage_170;
      dark_weights_normed_gauss_blur_3_update_0_stage_172 <= dark_weights_normed_gauss_blur_3_update_0_stage_171;
      dark_weights_normed_gauss_blur_3_update_0_stage_173 <= dark_weights_normed_gauss_blur_3_update_0_stage_172;
      dark_weights_normed_gauss_blur_3_update_0_stage_174 <= dark_weights_normed_gauss_blur_3_update_0_stage_173;
      dark_weights_normed_gauss_blur_3_update_0_stage_175 <= dark_weights_normed_gauss_blur_3_update_0_stage_174;
      dark_weights_normed_gauss_blur_3_update_0_stage_176 <= dark_weights_normed_gauss_blur_3_update_0_stage_175;
      dark_weights_normed_gauss_blur_3_update_0_stage_177 <= dark_weights_normed_gauss_blur_3_update_0_stage_176;
      dark_weights_normed_gauss_blur_3_update_0_stage_178 <= dark_weights_normed_gauss_blur_3_update_0_stage_177;
      dark_weights_normed_gauss_blur_3_update_0_stage_179 <= dark_weights_normed_gauss_blur_3_update_0_stage_178;
      dark_weights_normed_gauss_blur_3_update_0_stage_180 <= dark_weights_normed_gauss_blur_3_update_0_stage_179;
      dark_weights_normed_gauss_blur_3_update_0_stage_181 <= dark_weights_normed_gauss_blur_3_update_0_stage_180;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_109 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_110 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_109;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_111 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_110;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_112 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_111;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_113 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_112;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_114 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_113;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_115 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_114;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_116 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_115;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_117 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_116;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_118 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_117;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_119 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_118;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_120 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_119;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_121 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_120;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_122 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_121;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_123 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_122;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_124 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_123;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_125 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_124;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_126 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_125;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_127 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_126;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_128 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_127;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_129 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_128;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_130 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_129;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_131 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_130;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_132 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_131;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_133 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_132;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_134 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_133;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_135 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_134;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_136 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_135;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_137 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_136;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_138 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_137;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_139 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_138;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_140 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_139;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_141 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_140;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_142 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_141;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_143 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_142;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_144 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_143;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_145 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_144;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_146 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_145;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_147 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_146;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_148 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_147;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_149 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_148;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_150 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_149;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_151 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_150;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_152 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_151;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_153 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_152;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_154 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_153;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_155 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_154;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_156 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_155;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_157 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_156;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_158 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_157;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_159 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_158;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_160 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_159;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_161 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_160;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_162 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_161;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_163 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_162;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_164 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_163;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_165 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_164;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_166 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_165;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_167 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_166;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_168 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_167;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_169 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_168;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_170 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_169;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_171 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_170;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_172 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_171;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_173 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_172;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_174 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_173;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_175 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_174;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_176 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_175;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_177 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_176;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_178 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_177;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_179 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_178;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_180 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_179;
      dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_181 <= dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73_stage_180;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_110 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_111 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_110;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_112 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_111;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_113 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_112;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_114 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_113;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_115 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_114;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_116 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_115;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_117 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_116;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_118 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_117;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_119 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_118;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_120 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_119;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_121 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_120;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_122 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_121;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_123 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_122;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_124 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_123;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_125 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_124;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_126 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_125;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_127 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_126;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_128 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_127;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_129 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_128;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_130 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_129;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_131 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_130;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_132 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_131;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_133 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_132;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_134 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_133;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_135 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_134;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_136 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_135;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_137 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_136;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_138 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_137;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_139 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_138;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_140 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_139;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_141 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_140;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_142 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_141;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_143 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_142;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_144 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_143;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_145 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_144;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_146 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_145;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_147 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_146;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_148 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_147;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_149 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_148;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_150 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_149;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_151 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_150;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_152 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_151;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_153 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_152;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_154 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_153;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_155 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_154;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_156 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_155;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_157 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_156;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_158 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_157;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_159 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_158;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_160 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_159;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_161 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_160;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_162 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_161;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_163 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_162;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_164 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_163;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_165 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_164;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_166 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_165;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_167 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_166;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_168 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_167;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_169 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_168;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_170 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_169;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_171 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_170;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_172 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_171;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_173 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_172;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_174 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_173;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_175 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_174;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_176 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_175;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_177 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_176;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_178 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_177;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_179 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_178;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_180 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_179;
      dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_181 <= dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74_stage_180;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_111 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_112 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_111;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_113 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_112;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_114 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_113;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_115 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_114;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_116 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_115;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_117 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_116;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_118 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_117;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_119 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_118;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_120 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_119;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_121 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_120;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_122 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_121;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_123 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_122;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_124 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_123;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_125 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_124;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_126 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_125;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_127 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_126;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_128 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_127;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_129 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_128;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_130 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_129;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_131 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_130;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_132 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_131;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_133 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_132;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_134 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_133;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_135 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_134;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_136 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_135;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_137 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_136;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_138 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_137;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_139 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_138;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_140 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_139;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_141 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_140;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_142 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_141;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_143 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_142;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_144 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_143;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_145 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_144;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_146 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_145;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_147 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_146;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_148 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_147;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_149 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_148;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_150 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_149;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_151 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_150;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_152 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_151;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_153 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_152;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_154 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_153;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_155 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_154;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_156 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_155;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_157 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_156;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_158 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_157;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_159 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_158;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_160 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_159;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_161 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_160;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_162 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_161;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_163 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_162;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_164 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_163;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_165 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_164;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_166 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_165;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_167 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_166;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_168 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_167;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_169 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_168;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_170 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_169;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_171 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_170;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_172 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_171;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_173 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_172;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_174 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_173;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_175 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_174;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_176 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_175;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_177 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_176;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_178 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_177;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_179 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_178;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_180 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_179;
      dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_181 <= dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75_stage_180;
      dark_laplace_diff_1_update_0_stage_112 <= dark_laplace_diff_1_update_0;
      dark_laplace_diff_1_update_0_stage_113 <= dark_laplace_diff_1_update_0_stage_112;
      dark_laplace_diff_1_update_0_stage_114 <= dark_laplace_diff_1_update_0_stage_113;
      dark_laplace_diff_1_update_0_stage_115 <= dark_laplace_diff_1_update_0_stage_114;
      dark_laplace_diff_1_update_0_stage_116 <= dark_laplace_diff_1_update_0_stage_115;
      dark_laplace_diff_1_update_0_stage_117 <= dark_laplace_diff_1_update_0_stage_116;
      dark_laplace_diff_1_update_0_stage_118 <= dark_laplace_diff_1_update_0_stage_117;
      dark_laplace_diff_1_update_0_stage_119 <= dark_laplace_diff_1_update_0_stage_118;
      dark_laplace_diff_1_update_0_stage_120 <= dark_laplace_diff_1_update_0_stage_119;
      dark_laplace_diff_1_update_0_stage_121 <= dark_laplace_diff_1_update_0_stage_120;
      dark_laplace_diff_1_update_0_stage_122 <= dark_laplace_diff_1_update_0_stage_121;
      dark_laplace_diff_1_update_0_stage_123 <= dark_laplace_diff_1_update_0_stage_122;
      dark_laplace_diff_1_update_0_stage_124 <= dark_laplace_diff_1_update_0_stage_123;
      dark_laplace_diff_1_update_0_stage_125 <= dark_laplace_diff_1_update_0_stage_124;
      dark_laplace_diff_1_update_0_stage_126 <= dark_laplace_diff_1_update_0_stage_125;
      dark_laplace_diff_1_update_0_stage_127 <= dark_laplace_diff_1_update_0_stage_126;
      dark_laplace_diff_1_update_0_stage_128 <= dark_laplace_diff_1_update_0_stage_127;
      dark_laplace_diff_1_update_0_stage_129 <= dark_laplace_diff_1_update_0_stage_128;
      dark_laplace_diff_1_update_0_stage_130 <= dark_laplace_diff_1_update_0_stage_129;
      dark_laplace_diff_1_update_0_stage_131 <= dark_laplace_diff_1_update_0_stage_130;
      dark_laplace_diff_1_update_0_stage_132 <= dark_laplace_diff_1_update_0_stage_131;
      dark_laplace_diff_1_update_0_stage_133 <= dark_laplace_diff_1_update_0_stage_132;
      dark_laplace_diff_1_update_0_stage_134 <= dark_laplace_diff_1_update_0_stage_133;
      dark_laplace_diff_1_update_0_stage_135 <= dark_laplace_diff_1_update_0_stage_134;
      dark_laplace_diff_1_update_0_stage_136 <= dark_laplace_diff_1_update_0_stage_135;
      dark_laplace_diff_1_update_0_stage_137 <= dark_laplace_diff_1_update_0_stage_136;
      dark_laplace_diff_1_update_0_stage_138 <= dark_laplace_diff_1_update_0_stage_137;
      dark_laplace_diff_1_update_0_stage_139 <= dark_laplace_diff_1_update_0_stage_138;
      dark_laplace_diff_1_update_0_stage_140 <= dark_laplace_diff_1_update_0_stage_139;
      dark_laplace_diff_1_update_0_stage_141 <= dark_laplace_diff_1_update_0_stage_140;
      dark_laplace_diff_1_update_0_stage_142 <= dark_laplace_diff_1_update_0_stage_141;
      dark_laplace_diff_1_update_0_stage_143 <= dark_laplace_diff_1_update_0_stage_142;
      dark_laplace_diff_1_update_0_stage_144 <= dark_laplace_diff_1_update_0_stage_143;
      dark_laplace_diff_1_update_0_stage_145 <= dark_laplace_diff_1_update_0_stage_144;
      dark_laplace_diff_1_update_0_stage_146 <= dark_laplace_diff_1_update_0_stage_145;
      dark_laplace_diff_1_update_0_stage_147 <= dark_laplace_diff_1_update_0_stage_146;
      dark_laplace_diff_1_update_0_stage_148 <= dark_laplace_diff_1_update_0_stage_147;
      dark_laplace_diff_1_update_0_stage_149 <= dark_laplace_diff_1_update_0_stage_148;
      dark_laplace_diff_1_update_0_stage_150 <= dark_laplace_diff_1_update_0_stage_149;
      dark_laplace_diff_1_update_0_stage_151 <= dark_laplace_diff_1_update_0_stage_150;
      dark_laplace_diff_1_update_0_stage_152 <= dark_laplace_diff_1_update_0_stage_151;
      dark_laplace_diff_1_update_0_stage_153 <= dark_laplace_diff_1_update_0_stage_152;
      dark_laplace_diff_1_update_0_stage_154 <= dark_laplace_diff_1_update_0_stage_153;
      dark_laplace_diff_1_update_0_stage_155 <= dark_laplace_diff_1_update_0_stage_154;
      dark_laplace_diff_1_update_0_stage_156 <= dark_laplace_diff_1_update_0_stage_155;
      dark_laplace_diff_1_update_0_stage_157 <= dark_laplace_diff_1_update_0_stage_156;
      dark_laplace_diff_1_update_0_stage_158 <= dark_laplace_diff_1_update_0_stage_157;
      dark_laplace_diff_1_update_0_stage_159 <= dark_laplace_diff_1_update_0_stage_158;
      dark_laplace_diff_1_update_0_stage_160 <= dark_laplace_diff_1_update_0_stage_159;
      dark_laplace_diff_1_update_0_stage_161 <= dark_laplace_diff_1_update_0_stage_160;
      dark_laplace_diff_1_update_0_stage_162 <= dark_laplace_diff_1_update_0_stage_161;
      dark_laplace_diff_1_update_0_stage_163 <= dark_laplace_diff_1_update_0_stage_162;
      dark_laplace_diff_1_update_0_stage_164 <= dark_laplace_diff_1_update_0_stage_163;
      dark_laplace_diff_1_update_0_stage_165 <= dark_laplace_diff_1_update_0_stage_164;
      dark_laplace_diff_1_update_0_stage_166 <= dark_laplace_diff_1_update_0_stage_165;
      dark_laplace_diff_1_update_0_stage_167 <= dark_laplace_diff_1_update_0_stage_166;
      dark_laplace_diff_1_update_0_stage_168 <= dark_laplace_diff_1_update_0_stage_167;
      dark_laplace_diff_1_update_0_stage_169 <= dark_laplace_diff_1_update_0_stage_168;
      dark_laplace_diff_1_update_0_stage_170 <= dark_laplace_diff_1_update_0_stage_169;
      dark_laplace_diff_1_update_0_stage_171 <= dark_laplace_diff_1_update_0_stage_170;
      dark_laplace_diff_1_update_0_stage_172 <= dark_laplace_diff_1_update_0_stage_171;
      dark_laplace_diff_1_update_0_stage_173 <= dark_laplace_diff_1_update_0_stage_172;
      dark_laplace_diff_1_update_0_stage_174 <= dark_laplace_diff_1_update_0_stage_173;
      dark_laplace_diff_1_update_0_stage_175 <= dark_laplace_diff_1_update_0_stage_174;
      dark_laplace_diff_1_update_0_stage_176 <= dark_laplace_diff_1_update_0_stage_175;
      dark_laplace_diff_1_update_0_stage_177 <= dark_laplace_diff_1_update_0_stage_176;
      dark_laplace_diff_1_update_0_stage_178 <= dark_laplace_diff_1_update_0_stage_177;
      dark_laplace_diff_1_update_0_stage_179 <= dark_laplace_diff_1_update_0_stage_178;
      dark_laplace_diff_1_update_0_stage_180 <= dark_laplace_diff_1_update_0_stage_179;
      dark_laplace_diff_1_update_0_stage_181 <= dark_laplace_diff_1_update_0_stage_180;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_113 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_114 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_113;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_115 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_114;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_116 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_115;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_117 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_116;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_118 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_117;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_119 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_118;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_120 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_119;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_121 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_120;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_122 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_121;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_123 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_122;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_124 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_123;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_125 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_124;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_126 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_125;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_127 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_126;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_128 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_127;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_129 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_128;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_130 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_129;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_131 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_130;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_132 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_131;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_133 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_132;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_134 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_133;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_135 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_134;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_136 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_135;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_137 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_136;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_138 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_137;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_139 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_138;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_140 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_139;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_141 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_140;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_142 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_141;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_143 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_142;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_144 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_143;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_145 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_144;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_146 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_145;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_147 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_146;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_148 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_147;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_149 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_148;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_150 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_149;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_151 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_150;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_152 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_151;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_153 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_152;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_154 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_153;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_155 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_154;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_156 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_155;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_157 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_156;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_158 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_157;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_159 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_158;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_160 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_159;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_161 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_160;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_162 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_161;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_163 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_162;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_164 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_163;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_165 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_164;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_166 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_165;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_167 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_166;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_168 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_167;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_169 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_168;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_170 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_169;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_171 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_170;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_172 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_171;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_173 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_172;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_174 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_173;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_175 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_174;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_176 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_175;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_177 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_176;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_178 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_177;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_179 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_178;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_180 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_179;
      dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_181 <= dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76_stage_180;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_120 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_121 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_120;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_122 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_121;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_123 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_122;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_124 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_123;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_125 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_124;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_126 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_125;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_127 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_126;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_128 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_127;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_129 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_128;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_130 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_129;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_131 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_130;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_132 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_131;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_133 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_132;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_134 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_133;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_135 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_134;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_136 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_135;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_137 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_136;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_138 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_137;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_139 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_138;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_140 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_139;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_141 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_140;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_142 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_141;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_143 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_142;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_144 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_143;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_145 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_144;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_146 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_145;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_147 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_146;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_148 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_147;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_149 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_148;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_150 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_149;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_151 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_150;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_152 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_151;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_153 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_152;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_154 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_153;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_155 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_154;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_156 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_155;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_157 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_156;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_158 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_157;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_159 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_158;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_160 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_159;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_161 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_160;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_162 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_161;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_163 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_162;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_164 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_163;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_165 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_164;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_166 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_165;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_167 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_166;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_168 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_167;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_169 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_168;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_170 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_169;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_171 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_170;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_172 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_171;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_173 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_172;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_174 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_173;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_175 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_174;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_176 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_175;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_177 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_176;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_178 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_177;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_179 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_178;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_180 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_179;
      bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_181 <= bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82_stage_180;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_114 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_115 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_114;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_116 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_115;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_117 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_116;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_118 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_117;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_119 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_118;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_120 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_119;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_121 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_120;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_122 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_121;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_123 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_122;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_124 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_123;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_125 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_124;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_126 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_125;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_127 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_126;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_128 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_127;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_129 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_128;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_130 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_129;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_131 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_130;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_132 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_131;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_133 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_132;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_134 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_133;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_135 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_134;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_136 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_135;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_137 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_136;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_138 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_137;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_139 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_138;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_140 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_139;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_141 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_140;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_142 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_141;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_143 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_142;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_144 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_143;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_145 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_144;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_146 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_145;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_147 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_146;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_148 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_147;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_149 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_148;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_150 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_149;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_151 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_150;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_152 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_151;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_153 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_152;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_154 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_153;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_155 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_154;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_156 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_155;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_157 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_156;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_158 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_157;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_159 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_158;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_160 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_159;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_161 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_160;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_162 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_161;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_163 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_162;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_164 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_163;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_165 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_164;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_166 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_165;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_167 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_166;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_168 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_167;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_169 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_168;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_170 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_169;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_171 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_170;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_172 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_171;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_173 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_172;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_174 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_173;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_175 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_174;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_176 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_175;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_177 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_176;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_178 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_177;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_179 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_178;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_180 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_179;
      bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_181 <= bright_laplace_diff_0_fused_level_0_update_0_read_read_77_stage_180;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_115 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_116 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_115;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_117 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_116;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_118 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_117;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_119 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_118;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_120 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_119;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_121 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_120;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_122 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_121;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_123 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_122;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_124 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_123;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_125 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_124;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_126 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_125;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_127 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_126;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_128 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_127;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_129 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_128;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_130 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_129;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_131 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_130;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_132 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_131;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_133 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_132;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_134 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_133;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_135 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_134;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_136 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_135;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_137 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_136;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_138 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_137;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_139 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_138;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_140 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_139;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_141 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_140;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_142 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_141;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_143 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_142;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_144 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_143;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_145 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_144;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_146 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_145;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_147 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_146;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_148 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_147;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_149 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_148;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_150 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_149;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_151 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_150;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_152 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_151;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_153 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_152;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_154 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_153;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_155 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_154;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_156 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_155;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_157 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_156;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_158 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_157;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_159 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_158;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_160 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_159;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_161 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_160;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_162 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_161;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_163 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_162;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_164 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_163;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_165 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_164;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_166 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_165;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_167 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_166;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_168 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_167;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_169 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_168;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_170 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_169;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_171 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_170;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_172 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_171;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_173 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_172;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_174 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_173;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_175 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_174;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_176 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_175;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_177 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_176;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_178 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_177;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_179 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_178;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_180 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_179;
      dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_181 <= dark_laplace_diff_0_fused_level_0_update_0_read_read_78_stage_180;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_116 <= bright_weights_normed_fused_level_0_update_0_read_read_79;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_117 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_116;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_118 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_117;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_119 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_118;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_120 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_119;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_121 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_120;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_122 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_121;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_123 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_122;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_124 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_123;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_125 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_124;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_126 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_125;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_127 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_126;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_128 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_127;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_129 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_128;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_130 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_129;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_131 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_130;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_132 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_131;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_133 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_132;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_134 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_133;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_135 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_134;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_136 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_135;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_137 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_136;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_138 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_137;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_139 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_138;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_140 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_139;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_141 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_140;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_142 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_141;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_143 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_142;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_144 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_143;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_145 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_144;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_146 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_145;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_147 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_146;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_148 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_147;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_149 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_148;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_150 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_149;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_151 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_150;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_152 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_151;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_153 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_152;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_154 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_153;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_155 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_154;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_156 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_155;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_157 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_156;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_158 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_157;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_159 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_158;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_160 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_159;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_161 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_160;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_162 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_161;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_163 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_162;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_164 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_163;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_165 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_164;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_166 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_165;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_167 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_166;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_168 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_167;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_169 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_168;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_170 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_169;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_171 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_170;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_172 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_171;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_173 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_172;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_174 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_173;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_175 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_174;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_176 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_175;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_177 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_176;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_178 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_177;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_179 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_178;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_180 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_179;
      bright_weights_normed_fused_level_0_update_0_read_read_79_stage_181 <= bright_weights_normed_fused_level_0_update_0_read_read_79_stage_180;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_117 <= dark_weights_normed_fused_level_0_update_0_read_read_80;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_118 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_117;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_119 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_118;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_120 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_119;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_121 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_120;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_122 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_121;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_123 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_122;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_124 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_123;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_125 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_124;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_126 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_125;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_127 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_126;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_128 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_127;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_129 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_128;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_130 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_129;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_131 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_130;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_132 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_131;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_133 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_132;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_134 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_133;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_135 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_134;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_136 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_135;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_137 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_136;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_138 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_137;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_139 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_138;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_140 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_139;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_141 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_140;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_142 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_141;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_143 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_142;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_144 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_143;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_145 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_144;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_146 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_145;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_147 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_146;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_148 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_147;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_149 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_148;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_150 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_149;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_151 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_150;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_152 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_151;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_153 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_152;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_154 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_153;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_155 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_154;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_156 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_155;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_157 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_156;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_158 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_157;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_159 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_158;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_160 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_159;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_161 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_160;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_162 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_161;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_163 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_162;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_164 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_163;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_165 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_164;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_166 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_165;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_167 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_166;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_168 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_167;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_169 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_168;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_170 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_169;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_171 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_170;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_172 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_171;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_173 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_172;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_174 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_173;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_175 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_174;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_176 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_175;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_177 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_176;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_178 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_177;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_179 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_178;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_180 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_179;
      dark_weights_normed_fused_level_0_update_0_read_read_80_stage_181 <= dark_weights_normed_fused_level_0_update_0_read_read_80_stage_180;
      fused_level_0_update_0_stage_118 <= fused_level_0_update_0;
      fused_level_0_update_0_stage_119 <= fused_level_0_update_0_stage_118;
      fused_level_0_update_0_stage_120 <= fused_level_0_update_0_stage_119;
      fused_level_0_update_0_stage_121 <= fused_level_0_update_0_stage_120;
      fused_level_0_update_0_stage_122 <= fused_level_0_update_0_stage_121;
      fused_level_0_update_0_stage_123 <= fused_level_0_update_0_stage_122;
      fused_level_0_update_0_stage_124 <= fused_level_0_update_0_stage_123;
      fused_level_0_update_0_stage_125 <= fused_level_0_update_0_stage_124;
      fused_level_0_update_0_stage_126 <= fused_level_0_update_0_stage_125;
      fused_level_0_update_0_stage_127 <= fused_level_0_update_0_stage_126;
      fused_level_0_update_0_stage_128 <= fused_level_0_update_0_stage_127;
      fused_level_0_update_0_stage_129 <= fused_level_0_update_0_stage_128;
      fused_level_0_update_0_stage_130 <= fused_level_0_update_0_stage_129;
      fused_level_0_update_0_stage_131 <= fused_level_0_update_0_stage_130;
      fused_level_0_update_0_stage_132 <= fused_level_0_update_0_stage_131;
      fused_level_0_update_0_stage_133 <= fused_level_0_update_0_stage_132;
      fused_level_0_update_0_stage_134 <= fused_level_0_update_0_stage_133;
      fused_level_0_update_0_stage_135 <= fused_level_0_update_0_stage_134;
      fused_level_0_update_0_stage_136 <= fused_level_0_update_0_stage_135;
      fused_level_0_update_0_stage_137 <= fused_level_0_update_0_stage_136;
      fused_level_0_update_0_stage_138 <= fused_level_0_update_0_stage_137;
      fused_level_0_update_0_stage_139 <= fused_level_0_update_0_stage_138;
      fused_level_0_update_0_stage_140 <= fused_level_0_update_0_stage_139;
      fused_level_0_update_0_stage_141 <= fused_level_0_update_0_stage_140;
      fused_level_0_update_0_stage_142 <= fused_level_0_update_0_stage_141;
      fused_level_0_update_0_stage_143 <= fused_level_0_update_0_stage_142;
      fused_level_0_update_0_stage_144 <= fused_level_0_update_0_stage_143;
      fused_level_0_update_0_stage_145 <= fused_level_0_update_0_stage_144;
      fused_level_0_update_0_stage_146 <= fused_level_0_update_0_stage_145;
      fused_level_0_update_0_stage_147 <= fused_level_0_update_0_stage_146;
      fused_level_0_update_0_stage_148 <= fused_level_0_update_0_stage_147;
      fused_level_0_update_0_stage_149 <= fused_level_0_update_0_stage_148;
      fused_level_0_update_0_stage_150 <= fused_level_0_update_0_stage_149;
      fused_level_0_update_0_stage_151 <= fused_level_0_update_0_stage_150;
      fused_level_0_update_0_stage_152 <= fused_level_0_update_0_stage_151;
      fused_level_0_update_0_stage_153 <= fused_level_0_update_0_stage_152;
      fused_level_0_update_0_stage_154 <= fused_level_0_update_0_stage_153;
      fused_level_0_update_0_stage_155 <= fused_level_0_update_0_stage_154;
      fused_level_0_update_0_stage_156 <= fused_level_0_update_0_stage_155;
      fused_level_0_update_0_stage_157 <= fused_level_0_update_0_stage_156;
      fused_level_0_update_0_stage_158 <= fused_level_0_update_0_stage_157;
      fused_level_0_update_0_stage_159 <= fused_level_0_update_0_stage_158;
      fused_level_0_update_0_stage_160 <= fused_level_0_update_0_stage_159;
      fused_level_0_update_0_stage_161 <= fused_level_0_update_0_stage_160;
      fused_level_0_update_0_stage_162 <= fused_level_0_update_0_stage_161;
      fused_level_0_update_0_stage_163 <= fused_level_0_update_0_stage_162;
      fused_level_0_update_0_stage_164 <= fused_level_0_update_0_stage_163;
      fused_level_0_update_0_stage_165 <= fused_level_0_update_0_stage_164;
      fused_level_0_update_0_stage_166 <= fused_level_0_update_0_stage_165;
      fused_level_0_update_0_stage_167 <= fused_level_0_update_0_stage_166;
      fused_level_0_update_0_stage_168 <= fused_level_0_update_0_stage_167;
      fused_level_0_update_0_stage_169 <= fused_level_0_update_0_stage_168;
      fused_level_0_update_0_stage_170 <= fused_level_0_update_0_stage_169;
      fused_level_0_update_0_stage_171 <= fused_level_0_update_0_stage_170;
      fused_level_0_update_0_stage_172 <= fused_level_0_update_0_stage_171;
      fused_level_0_update_0_stage_173 <= fused_level_0_update_0_stage_172;
      fused_level_0_update_0_stage_174 <= fused_level_0_update_0_stage_173;
      fused_level_0_update_0_stage_175 <= fused_level_0_update_0_stage_174;
      fused_level_0_update_0_stage_176 <= fused_level_0_update_0_stage_175;
      fused_level_0_update_0_stage_177 <= fused_level_0_update_0_stage_176;
      fused_level_0_update_0_stage_178 <= fused_level_0_update_0_stage_177;
      fused_level_0_update_0_stage_179 <= fused_level_0_update_0_stage_178;
      fused_level_0_update_0_stage_180 <= fused_level_0_update_0_stage_179;
      fused_level_0_update_0_stage_181 <= fused_level_0_update_0_stage_180;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_119 <= fused_level_0_fused_level_0_update_0_write_write_81;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_120 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_119;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_121 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_120;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_122 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_121;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_123 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_122;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_124 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_123;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_125 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_124;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_126 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_125;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_127 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_126;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_128 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_127;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_129 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_128;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_130 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_129;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_131 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_130;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_132 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_131;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_133 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_132;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_134 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_133;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_135 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_134;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_136 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_135;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_137 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_136;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_138 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_137;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_139 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_138;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_140 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_139;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_141 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_140;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_142 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_141;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_143 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_142;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_144 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_143;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_145 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_144;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_146 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_145;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_147 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_146;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_148 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_147;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_149 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_148;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_150 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_149;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_151 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_150;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_152 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_151;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_153 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_152;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_154 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_153;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_155 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_154;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_156 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_155;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_157 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_156;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_158 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_157;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_159 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_158;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_160 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_159;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_161 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_160;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_162 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_161;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_163 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_162;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_164 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_163;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_165 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_164;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_166 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_165;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_167 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_166;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_168 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_167;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_169 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_168;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_170 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_169;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_171 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_170;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_172 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_171;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_173 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_172;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_174 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_173;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_175 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_174;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_176 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_175;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_177 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_176;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_178 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_177;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_179 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_178;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_180 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_179;
      fused_level_0_fused_level_0_update_0_write_write_81_stage_181 <= fused_level_0_fused_level_0_update_0_write_write_81_stage_180;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_121 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_122 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_121;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_123 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_122;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_124 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_123;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_125 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_124;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_126 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_125;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_127 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_126;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_128 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_127;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_129 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_128;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_130 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_129;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_131 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_130;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_132 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_131;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_133 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_132;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_134 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_133;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_135 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_134;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_136 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_135;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_137 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_136;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_138 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_137;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_139 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_138;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_140 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_139;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_141 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_140;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_142 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_141;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_143 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_142;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_144 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_143;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_145 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_144;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_146 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_145;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_147 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_146;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_148 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_147;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_149 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_148;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_150 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_149;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_151 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_150;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_152 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_151;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_153 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_152;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_154 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_153;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_155 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_154;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_156 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_155;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_157 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_156;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_158 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_157;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_159 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_158;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_160 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_159;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_161 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_160;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_162 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_161;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_163 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_162;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_164 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_163;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_165 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_164;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_166 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_165;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_167 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_166;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_168 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_167;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_169 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_168;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_170 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_169;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_171 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_170;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_172 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_171;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_173 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_172;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_174 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_173;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_175 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_174;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_176 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_175;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_177 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_176;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_178 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_177;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_179 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_178;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_180 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_179;
      bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_181 <= bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83_stage_180;
      bright_laplace_diff_2_update_0_stage_122 <= bright_laplace_diff_2_update_0;
      bright_laplace_diff_2_update_0_stage_123 <= bright_laplace_diff_2_update_0_stage_122;
      bright_laplace_diff_2_update_0_stage_124 <= bright_laplace_diff_2_update_0_stage_123;
      bright_laplace_diff_2_update_0_stage_125 <= bright_laplace_diff_2_update_0_stage_124;
      bright_laplace_diff_2_update_0_stage_126 <= bright_laplace_diff_2_update_0_stage_125;
      bright_laplace_diff_2_update_0_stage_127 <= bright_laplace_diff_2_update_0_stage_126;
      bright_laplace_diff_2_update_0_stage_128 <= bright_laplace_diff_2_update_0_stage_127;
      bright_laplace_diff_2_update_0_stage_129 <= bright_laplace_diff_2_update_0_stage_128;
      bright_laplace_diff_2_update_0_stage_130 <= bright_laplace_diff_2_update_0_stage_129;
      bright_laplace_diff_2_update_0_stage_131 <= bright_laplace_diff_2_update_0_stage_130;
      bright_laplace_diff_2_update_0_stage_132 <= bright_laplace_diff_2_update_0_stage_131;
      bright_laplace_diff_2_update_0_stage_133 <= bright_laplace_diff_2_update_0_stage_132;
      bright_laplace_diff_2_update_0_stage_134 <= bright_laplace_diff_2_update_0_stage_133;
      bright_laplace_diff_2_update_0_stage_135 <= bright_laplace_diff_2_update_0_stage_134;
      bright_laplace_diff_2_update_0_stage_136 <= bright_laplace_diff_2_update_0_stage_135;
      bright_laplace_diff_2_update_0_stage_137 <= bright_laplace_diff_2_update_0_stage_136;
      bright_laplace_diff_2_update_0_stage_138 <= bright_laplace_diff_2_update_0_stage_137;
      bright_laplace_diff_2_update_0_stage_139 <= bright_laplace_diff_2_update_0_stage_138;
      bright_laplace_diff_2_update_0_stage_140 <= bright_laplace_diff_2_update_0_stage_139;
      bright_laplace_diff_2_update_0_stage_141 <= bright_laplace_diff_2_update_0_stage_140;
      bright_laplace_diff_2_update_0_stage_142 <= bright_laplace_diff_2_update_0_stage_141;
      bright_laplace_diff_2_update_0_stage_143 <= bright_laplace_diff_2_update_0_stage_142;
      bright_laplace_diff_2_update_0_stage_144 <= bright_laplace_diff_2_update_0_stage_143;
      bright_laplace_diff_2_update_0_stage_145 <= bright_laplace_diff_2_update_0_stage_144;
      bright_laplace_diff_2_update_0_stage_146 <= bright_laplace_diff_2_update_0_stage_145;
      bright_laplace_diff_2_update_0_stage_147 <= bright_laplace_diff_2_update_0_stage_146;
      bright_laplace_diff_2_update_0_stage_148 <= bright_laplace_diff_2_update_0_stage_147;
      bright_laplace_diff_2_update_0_stage_149 <= bright_laplace_diff_2_update_0_stage_148;
      bright_laplace_diff_2_update_0_stage_150 <= bright_laplace_diff_2_update_0_stage_149;
      bright_laplace_diff_2_update_0_stage_151 <= bright_laplace_diff_2_update_0_stage_150;
      bright_laplace_diff_2_update_0_stage_152 <= bright_laplace_diff_2_update_0_stage_151;
      bright_laplace_diff_2_update_0_stage_153 <= bright_laplace_diff_2_update_0_stage_152;
      bright_laplace_diff_2_update_0_stage_154 <= bright_laplace_diff_2_update_0_stage_153;
      bright_laplace_diff_2_update_0_stage_155 <= bright_laplace_diff_2_update_0_stage_154;
      bright_laplace_diff_2_update_0_stage_156 <= bright_laplace_diff_2_update_0_stage_155;
      bright_laplace_diff_2_update_0_stage_157 <= bright_laplace_diff_2_update_0_stage_156;
      bright_laplace_diff_2_update_0_stage_158 <= bright_laplace_diff_2_update_0_stage_157;
      bright_laplace_diff_2_update_0_stage_159 <= bright_laplace_diff_2_update_0_stage_158;
      bright_laplace_diff_2_update_0_stage_160 <= bright_laplace_diff_2_update_0_stage_159;
      bright_laplace_diff_2_update_0_stage_161 <= bright_laplace_diff_2_update_0_stage_160;
      bright_laplace_diff_2_update_0_stage_162 <= bright_laplace_diff_2_update_0_stage_161;
      bright_laplace_diff_2_update_0_stage_163 <= bright_laplace_diff_2_update_0_stage_162;
      bright_laplace_diff_2_update_0_stage_164 <= bright_laplace_diff_2_update_0_stage_163;
      bright_laplace_diff_2_update_0_stage_165 <= bright_laplace_diff_2_update_0_stage_164;
      bright_laplace_diff_2_update_0_stage_166 <= bright_laplace_diff_2_update_0_stage_165;
      bright_laplace_diff_2_update_0_stage_167 <= bright_laplace_diff_2_update_0_stage_166;
      bright_laplace_diff_2_update_0_stage_168 <= bright_laplace_diff_2_update_0_stage_167;
      bright_laplace_diff_2_update_0_stage_169 <= bright_laplace_diff_2_update_0_stage_168;
      bright_laplace_diff_2_update_0_stage_170 <= bright_laplace_diff_2_update_0_stage_169;
      bright_laplace_diff_2_update_0_stage_171 <= bright_laplace_diff_2_update_0_stage_170;
      bright_laplace_diff_2_update_0_stage_172 <= bright_laplace_diff_2_update_0_stage_171;
      bright_laplace_diff_2_update_0_stage_173 <= bright_laplace_diff_2_update_0_stage_172;
      bright_laplace_diff_2_update_0_stage_174 <= bright_laplace_diff_2_update_0_stage_173;
      bright_laplace_diff_2_update_0_stage_175 <= bright_laplace_diff_2_update_0_stage_174;
      bright_laplace_diff_2_update_0_stage_176 <= bright_laplace_diff_2_update_0_stage_175;
      bright_laplace_diff_2_update_0_stage_177 <= bright_laplace_diff_2_update_0_stage_176;
      bright_laplace_diff_2_update_0_stage_178 <= bright_laplace_diff_2_update_0_stage_177;
      bright_laplace_diff_2_update_0_stage_179 <= bright_laplace_diff_2_update_0_stage_178;
      bright_laplace_diff_2_update_0_stage_180 <= bright_laplace_diff_2_update_0_stage_179;
      bright_laplace_diff_2_update_0_stage_181 <= bright_laplace_diff_2_update_0_stage_180;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_123 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_124 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_123;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_125 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_124;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_126 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_125;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_127 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_126;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_128 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_127;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_129 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_128;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_130 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_129;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_131 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_130;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_132 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_131;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_133 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_132;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_134 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_133;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_135 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_134;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_136 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_135;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_137 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_136;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_138 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_137;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_139 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_138;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_140 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_139;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_141 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_140;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_142 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_141;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_143 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_142;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_144 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_143;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_145 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_144;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_146 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_145;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_147 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_146;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_148 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_147;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_149 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_148;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_150 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_149;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_151 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_150;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_152 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_151;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_153 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_152;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_154 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_153;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_155 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_154;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_156 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_155;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_157 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_156;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_158 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_157;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_159 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_158;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_160 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_159;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_161 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_160;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_162 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_161;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_163 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_162;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_164 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_163;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_165 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_164;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_166 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_165;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_167 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_166;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_168 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_167;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_169 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_168;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_170 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_169;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_171 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_170;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_172 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_171;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_173 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_172;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_174 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_173;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_175 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_174;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_176 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_175;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_177 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_176;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_178 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_177;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_179 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_178;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_180 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_179;
      bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_181 <= bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84_stage_180;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_130 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_131 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_130;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_132 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_131;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_133 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_132;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_134 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_133;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_135 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_134;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_136 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_135;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_137 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_136;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_138 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_137;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_139 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_138;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_140 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_139;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_141 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_140;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_142 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_141;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_143 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_142;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_144 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_143;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_145 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_144;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_146 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_145;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_147 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_146;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_148 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_147;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_149 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_148;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_150 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_149;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_151 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_150;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_152 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_151;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_153 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_152;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_154 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_153;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_155 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_154;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_156 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_155;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_157 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_156;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_158 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_157;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_159 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_158;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_160 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_159;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_161 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_160;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_162 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_161;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_163 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_162;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_164 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_163;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_165 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_164;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_166 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_165;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_167 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_166;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_168 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_167;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_169 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_168;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_170 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_169;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_171 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_170;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_172 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_171;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_173 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_172;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_174 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_173;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_175 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_174;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_176 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_175;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_177 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_176;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_178 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_177;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_179 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_178;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_180 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_179;
      bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_181 <= bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90_stage_180;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_124 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_125 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_124;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_126 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_125;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_127 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_126;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_128 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_127;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_129 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_128;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_130 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_129;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_131 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_130;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_132 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_131;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_133 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_132;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_134 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_133;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_135 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_134;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_136 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_135;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_137 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_136;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_138 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_137;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_139 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_138;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_140 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_139;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_141 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_140;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_142 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_141;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_143 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_142;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_144 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_143;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_145 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_144;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_146 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_145;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_147 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_146;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_148 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_147;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_149 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_148;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_150 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_149;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_151 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_150;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_152 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_151;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_153 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_152;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_154 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_153;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_155 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_154;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_156 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_155;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_157 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_156;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_158 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_157;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_159 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_158;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_160 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_159;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_161 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_160;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_162 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_161;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_163 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_162;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_164 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_163;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_165 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_164;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_166 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_165;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_167 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_166;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_168 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_167;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_169 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_168;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_170 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_169;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_171 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_170;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_172 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_171;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_173 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_172;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_174 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_173;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_175 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_174;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_176 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_175;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_177 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_176;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_178 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_177;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_179 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_178;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_180 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_179;
      bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_181 <= bright_laplace_diff_1_fused_level_1_update_0_read_read_85_stage_180;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_125 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_126 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_125;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_127 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_126;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_128 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_127;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_129 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_128;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_130 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_129;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_131 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_130;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_132 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_131;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_133 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_132;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_134 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_133;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_135 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_134;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_136 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_135;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_137 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_136;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_138 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_137;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_139 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_138;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_140 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_139;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_141 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_140;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_142 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_141;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_143 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_142;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_144 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_143;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_145 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_144;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_146 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_145;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_147 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_146;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_148 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_147;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_149 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_148;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_150 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_149;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_151 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_150;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_152 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_151;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_153 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_152;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_154 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_153;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_155 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_154;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_156 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_155;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_157 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_156;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_158 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_157;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_159 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_158;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_160 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_159;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_161 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_160;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_162 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_161;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_163 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_162;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_164 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_163;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_165 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_164;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_166 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_165;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_167 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_166;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_168 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_167;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_169 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_168;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_170 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_169;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_171 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_170;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_172 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_171;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_173 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_172;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_174 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_173;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_175 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_174;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_176 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_175;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_177 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_176;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_178 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_177;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_179 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_178;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_180 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_179;
      dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_181 <= dark_laplace_diff_1_fused_level_1_update_0_read_read_86_stage_180;
      bright_weights_normed_gauss_blur_2_update_0_stage_131 <= bright_weights_normed_gauss_blur_2_update_0;
      bright_weights_normed_gauss_blur_2_update_0_stage_132 <= bright_weights_normed_gauss_blur_2_update_0_stage_131;
      bright_weights_normed_gauss_blur_2_update_0_stage_133 <= bright_weights_normed_gauss_blur_2_update_0_stage_132;
      bright_weights_normed_gauss_blur_2_update_0_stage_134 <= bright_weights_normed_gauss_blur_2_update_0_stage_133;
      bright_weights_normed_gauss_blur_2_update_0_stage_135 <= bright_weights_normed_gauss_blur_2_update_0_stage_134;
      bright_weights_normed_gauss_blur_2_update_0_stage_136 <= bright_weights_normed_gauss_blur_2_update_0_stage_135;
      bright_weights_normed_gauss_blur_2_update_0_stage_137 <= bright_weights_normed_gauss_blur_2_update_0_stage_136;
      bright_weights_normed_gauss_blur_2_update_0_stage_138 <= bright_weights_normed_gauss_blur_2_update_0_stage_137;
      bright_weights_normed_gauss_blur_2_update_0_stage_139 <= bright_weights_normed_gauss_blur_2_update_0_stage_138;
      bright_weights_normed_gauss_blur_2_update_0_stage_140 <= bright_weights_normed_gauss_blur_2_update_0_stage_139;
      bright_weights_normed_gauss_blur_2_update_0_stage_141 <= bright_weights_normed_gauss_blur_2_update_0_stage_140;
      bright_weights_normed_gauss_blur_2_update_0_stage_142 <= bright_weights_normed_gauss_blur_2_update_0_stage_141;
      bright_weights_normed_gauss_blur_2_update_0_stage_143 <= bright_weights_normed_gauss_blur_2_update_0_stage_142;
      bright_weights_normed_gauss_blur_2_update_0_stage_144 <= bright_weights_normed_gauss_blur_2_update_0_stage_143;
      bright_weights_normed_gauss_blur_2_update_0_stage_145 <= bright_weights_normed_gauss_blur_2_update_0_stage_144;
      bright_weights_normed_gauss_blur_2_update_0_stage_146 <= bright_weights_normed_gauss_blur_2_update_0_stage_145;
      bright_weights_normed_gauss_blur_2_update_0_stage_147 <= bright_weights_normed_gauss_blur_2_update_0_stage_146;
      bright_weights_normed_gauss_blur_2_update_0_stage_148 <= bright_weights_normed_gauss_blur_2_update_0_stage_147;
      bright_weights_normed_gauss_blur_2_update_0_stage_149 <= bright_weights_normed_gauss_blur_2_update_0_stage_148;
      bright_weights_normed_gauss_blur_2_update_0_stage_150 <= bright_weights_normed_gauss_blur_2_update_0_stage_149;
      bright_weights_normed_gauss_blur_2_update_0_stage_151 <= bright_weights_normed_gauss_blur_2_update_0_stage_150;
      bright_weights_normed_gauss_blur_2_update_0_stage_152 <= bright_weights_normed_gauss_blur_2_update_0_stage_151;
      bright_weights_normed_gauss_blur_2_update_0_stage_153 <= bright_weights_normed_gauss_blur_2_update_0_stage_152;
      bright_weights_normed_gauss_blur_2_update_0_stage_154 <= bright_weights_normed_gauss_blur_2_update_0_stage_153;
      bright_weights_normed_gauss_blur_2_update_0_stage_155 <= bright_weights_normed_gauss_blur_2_update_0_stage_154;
      bright_weights_normed_gauss_blur_2_update_0_stage_156 <= bright_weights_normed_gauss_blur_2_update_0_stage_155;
      bright_weights_normed_gauss_blur_2_update_0_stage_157 <= bright_weights_normed_gauss_blur_2_update_0_stage_156;
      bright_weights_normed_gauss_blur_2_update_0_stage_158 <= bright_weights_normed_gauss_blur_2_update_0_stage_157;
      bright_weights_normed_gauss_blur_2_update_0_stage_159 <= bright_weights_normed_gauss_blur_2_update_0_stage_158;
      bright_weights_normed_gauss_blur_2_update_0_stage_160 <= bright_weights_normed_gauss_blur_2_update_0_stage_159;
      bright_weights_normed_gauss_blur_2_update_0_stage_161 <= bright_weights_normed_gauss_blur_2_update_0_stage_160;
      bright_weights_normed_gauss_blur_2_update_0_stage_162 <= bright_weights_normed_gauss_blur_2_update_0_stage_161;
      bright_weights_normed_gauss_blur_2_update_0_stage_163 <= bright_weights_normed_gauss_blur_2_update_0_stage_162;
      bright_weights_normed_gauss_blur_2_update_0_stage_164 <= bright_weights_normed_gauss_blur_2_update_0_stage_163;
      bright_weights_normed_gauss_blur_2_update_0_stage_165 <= bright_weights_normed_gauss_blur_2_update_0_stage_164;
      bright_weights_normed_gauss_blur_2_update_0_stage_166 <= bright_weights_normed_gauss_blur_2_update_0_stage_165;
      bright_weights_normed_gauss_blur_2_update_0_stage_167 <= bright_weights_normed_gauss_blur_2_update_0_stage_166;
      bright_weights_normed_gauss_blur_2_update_0_stage_168 <= bright_weights_normed_gauss_blur_2_update_0_stage_167;
      bright_weights_normed_gauss_blur_2_update_0_stage_169 <= bright_weights_normed_gauss_blur_2_update_0_stage_168;
      bright_weights_normed_gauss_blur_2_update_0_stage_170 <= bright_weights_normed_gauss_blur_2_update_0_stage_169;
      bright_weights_normed_gauss_blur_2_update_0_stage_171 <= bright_weights_normed_gauss_blur_2_update_0_stage_170;
      bright_weights_normed_gauss_blur_2_update_0_stage_172 <= bright_weights_normed_gauss_blur_2_update_0_stage_171;
      bright_weights_normed_gauss_blur_2_update_0_stage_173 <= bright_weights_normed_gauss_blur_2_update_0_stage_172;
      bright_weights_normed_gauss_blur_2_update_0_stage_174 <= bright_weights_normed_gauss_blur_2_update_0_stage_173;
      bright_weights_normed_gauss_blur_2_update_0_stage_175 <= bright_weights_normed_gauss_blur_2_update_0_stage_174;
      bright_weights_normed_gauss_blur_2_update_0_stage_176 <= bright_weights_normed_gauss_blur_2_update_0_stage_175;
      bright_weights_normed_gauss_blur_2_update_0_stage_177 <= bright_weights_normed_gauss_blur_2_update_0_stage_176;
      bright_weights_normed_gauss_blur_2_update_0_stage_178 <= bright_weights_normed_gauss_blur_2_update_0_stage_177;
      bright_weights_normed_gauss_blur_2_update_0_stage_179 <= bright_weights_normed_gauss_blur_2_update_0_stage_178;
      bright_weights_normed_gauss_blur_2_update_0_stage_180 <= bright_weights_normed_gauss_blur_2_update_0_stage_179;
      bright_weights_normed_gauss_blur_2_update_0_stage_181 <= bright_weights_normed_gauss_blur_2_update_0_stage_180;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_133 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_134 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_133;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_135 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_134;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_136 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_135;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_137 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_136;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_138 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_137;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_139 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_138;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_140 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_139;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_141 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_140;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_142 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_141;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_143 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_142;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_144 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_143;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_145 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_144;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_146 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_145;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_147 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_146;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_148 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_147;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_149 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_148;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_150 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_149;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_151 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_150;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_152 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_151;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_153 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_152;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_154 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_153;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_155 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_154;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_156 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_155;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_157 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_156;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_158 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_157;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_159 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_158;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_160 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_159;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_161 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_160;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_162 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_161;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_163 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_162;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_164 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_163;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_165 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_164;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_166 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_165;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_167 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_166;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_168 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_167;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_169 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_168;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_170 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_169;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_171 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_170;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_172 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_171;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_173 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_172;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_174 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_173;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_175 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_174;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_176 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_175;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_177 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_176;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_178 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_177;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_179 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_178;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_180 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_179;
      dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_181 <= dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92_stage_180;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_132 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_133 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_132;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_134 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_133;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_135 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_134;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_136 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_135;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_137 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_136;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_138 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_137;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_139 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_138;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_140 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_139;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_141 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_140;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_142 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_141;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_143 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_142;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_144 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_143;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_145 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_144;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_146 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_145;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_147 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_146;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_148 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_147;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_149 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_148;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_150 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_149;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_151 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_150;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_152 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_151;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_153 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_152;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_154 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_153;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_155 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_154;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_156 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_155;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_157 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_156;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_158 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_157;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_159 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_158;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_160 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_159;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_161 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_160;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_162 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_161;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_163 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_162;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_164 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_163;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_165 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_164;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_166 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_165;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_167 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_166;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_168 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_167;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_169 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_168;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_170 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_169;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_171 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_170;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_172 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_171;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_173 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_172;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_174 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_173;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_175 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_174;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_176 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_175;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_177 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_176;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_178 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_177;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_179 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_178;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_180 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_179;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_181 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91_stage_180;
      dark_gauss_ds_3_update_0_stage_134 <= dark_gauss_ds_3_update_0;
      dark_gauss_ds_3_update_0_stage_135 <= dark_gauss_ds_3_update_0_stage_134;
      dark_gauss_ds_3_update_0_stage_136 <= dark_gauss_ds_3_update_0_stage_135;
      dark_gauss_ds_3_update_0_stage_137 <= dark_gauss_ds_3_update_0_stage_136;
      dark_gauss_ds_3_update_0_stage_138 <= dark_gauss_ds_3_update_0_stage_137;
      dark_gauss_ds_3_update_0_stage_139 <= dark_gauss_ds_3_update_0_stage_138;
      dark_gauss_ds_3_update_0_stage_140 <= dark_gauss_ds_3_update_0_stage_139;
      dark_gauss_ds_3_update_0_stage_141 <= dark_gauss_ds_3_update_0_stage_140;
      dark_gauss_ds_3_update_0_stage_142 <= dark_gauss_ds_3_update_0_stage_141;
      dark_gauss_ds_3_update_0_stage_143 <= dark_gauss_ds_3_update_0_stage_142;
      dark_gauss_ds_3_update_0_stage_144 <= dark_gauss_ds_3_update_0_stage_143;
      dark_gauss_ds_3_update_0_stage_145 <= dark_gauss_ds_3_update_0_stage_144;
      dark_gauss_ds_3_update_0_stage_146 <= dark_gauss_ds_3_update_0_stage_145;
      dark_gauss_ds_3_update_0_stage_147 <= dark_gauss_ds_3_update_0_stage_146;
      dark_gauss_ds_3_update_0_stage_148 <= dark_gauss_ds_3_update_0_stage_147;
      dark_gauss_ds_3_update_0_stage_149 <= dark_gauss_ds_3_update_0_stage_148;
      dark_gauss_ds_3_update_0_stage_150 <= dark_gauss_ds_3_update_0_stage_149;
      dark_gauss_ds_3_update_0_stage_151 <= dark_gauss_ds_3_update_0_stage_150;
      dark_gauss_ds_3_update_0_stage_152 <= dark_gauss_ds_3_update_0_stage_151;
      dark_gauss_ds_3_update_0_stage_153 <= dark_gauss_ds_3_update_0_stage_152;
      dark_gauss_ds_3_update_0_stage_154 <= dark_gauss_ds_3_update_0_stage_153;
      dark_gauss_ds_3_update_0_stage_155 <= dark_gauss_ds_3_update_0_stage_154;
      dark_gauss_ds_3_update_0_stage_156 <= dark_gauss_ds_3_update_0_stage_155;
      dark_gauss_ds_3_update_0_stage_157 <= dark_gauss_ds_3_update_0_stage_156;
      dark_gauss_ds_3_update_0_stage_158 <= dark_gauss_ds_3_update_0_stage_157;
      dark_gauss_ds_3_update_0_stage_159 <= dark_gauss_ds_3_update_0_stage_158;
      dark_gauss_ds_3_update_0_stage_160 <= dark_gauss_ds_3_update_0_stage_159;
      dark_gauss_ds_3_update_0_stage_161 <= dark_gauss_ds_3_update_0_stage_160;
      dark_gauss_ds_3_update_0_stage_162 <= dark_gauss_ds_3_update_0_stage_161;
      dark_gauss_ds_3_update_0_stage_163 <= dark_gauss_ds_3_update_0_stage_162;
      dark_gauss_ds_3_update_0_stage_164 <= dark_gauss_ds_3_update_0_stage_163;
      dark_gauss_ds_3_update_0_stage_165 <= dark_gauss_ds_3_update_0_stage_164;
      dark_gauss_ds_3_update_0_stage_166 <= dark_gauss_ds_3_update_0_stage_165;
      dark_gauss_ds_3_update_0_stage_167 <= dark_gauss_ds_3_update_0_stage_166;
      dark_gauss_ds_3_update_0_stage_168 <= dark_gauss_ds_3_update_0_stage_167;
      dark_gauss_ds_3_update_0_stage_169 <= dark_gauss_ds_3_update_0_stage_168;
      dark_gauss_ds_3_update_0_stage_170 <= dark_gauss_ds_3_update_0_stage_169;
      dark_gauss_ds_3_update_0_stage_171 <= dark_gauss_ds_3_update_0_stage_170;
      dark_gauss_ds_3_update_0_stage_172 <= dark_gauss_ds_3_update_0_stage_171;
      dark_gauss_ds_3_update_0_stage_173 <= dark_gauss_ds_3_update_0_stage_172;
      dark_gauss_ds_3_update_0_stage_174 <= dark_gauss_ds_3_update_0_stage_173;
      dark_gauss_ds_3_update_0_stage_175 <= dark_gauss_ds_3_update_0_stage_174;
      dark_gauss_ds_3_update_0_stage_176 <= dark_gauss_ds_3_update_0_stage_175;
      dark_gauss_ds_3_update_0_stage_177 <= dark_gauss_ds_3_update_0_stage_176;
      dark_gauss_ds_3_update_0_stage_178 <= dark_gauss_ds_3_update_0_stage_177;
      dark_gauss_ds_3_update_0_stage_179 <= dark_gauss_ds_3_update_0_stage_178;
      dark_gauss_ds_3_update_0_stage_180 <= dark_gauss_ds_3_update_0_stage_179;
      dark_gauss_ds_3_update_0_stage_181 <= dark_gauss_ds_3_update_0_stage_180;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_135 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_136 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_135;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_137 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_136;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_138 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_137;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_139 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_138;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_140 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_139;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_141 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_140;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_142 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_141;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_143 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_142;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_144 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_143;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_145 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_144;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_146 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_145;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_147 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_146;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_148 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_147;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_149 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_148;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_150 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_149;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_151 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_150;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_152 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_151;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_153 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_152;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_154 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_153;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_155 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_154;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_156 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_155;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_157 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_156;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_158 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_157;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_159 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_158;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_160 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_159;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_161 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_160;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_162 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_161;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_163 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_162;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_164 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_163;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_165 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_164;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_166 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_165;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_167 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_166;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_168 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_167;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_169 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_168;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_170 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_169;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_171 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_170;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_172 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_171;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_173 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_172;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_174 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_173;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_175 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_174;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_176 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_175;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_177 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_176;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_178 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_177;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_179 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_178;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_180 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_179;
      dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_181 <= dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93_stage_180;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_139 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_140 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_139;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_141 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_140;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_142 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_141;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_143 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_142;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_144 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_143;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_145 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_144;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_146 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_145;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_147 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_146;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_148 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_147;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_149 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_148;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_150 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_149;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_151 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_150;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_152 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_151;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_153 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_152;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_154 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_153;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_155 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_154;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_156 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_155;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_157 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_156;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_158 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_157;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_159 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_158;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_160 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_159;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_161 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_160;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_162 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_161;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_163 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_162;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_164 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_163;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_165 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_164;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_166 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_165;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_167 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_166;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_168 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_167;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_169 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_168;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_170 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_169;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_171 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_170;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_172 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_171;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_173 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_172;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_174 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_173;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_175 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_174;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_176 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_175;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_177 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_176;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_178 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_177;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_179 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_178;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_180 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_179;
      bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_181 <= bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96_stage_180;
      bright_weights_normed_gauss_ds_2_update_0_stage_140 <= bright_weights_normed_gauss_ds_2_update_0;
      bright_weights_normed_gauss_ds_2_update_0_stage_141 <= bright_weights_normed_gauss_ds_2_update_0_stage_140;
      bright_weights_normed_gauss_ds_2_update_0_stage_142 <= bright_weights_normed_gauss_ds_2_update_0_stage_141;
      bright_weights_normed_gauss_ds_2_update_0_stage_143 <= bright_weights_normed_gauss_ds_2_update_0_stage_142;
      bright_weights_normed_gauss_ds_2_update_0_stage_144 <= bright_weights_normed_gauss_ds_2_update_0_stage_143;
      bright_weights_normed_gauss_ds_2_update_0_stage_145 <= bright_weights_normed_gauss_ds_2_update_0_stage_144;
      bright_weights_normed_gauss_ds_2_update_0_stage_146 <= bright_weights_normed_gauss_ds_2_update_0_stage_145;
      bright_weights_normed_gauss_ds_2_update_0_stage_147 <= bright_weights_normed_gauss_ds_2_update_0_stage_146;
      bright_weights_normed_gauss_ds_2_update_0_stage_148 <= bright_weights_normed_gauss_ds_2_update_0_stage_147;
      bright_weights_normed_gauss_ds_2_update_0_stage_149 <= bright_weights_normed_gauss_ds_2_update_0_stage_148;
      bright_weights_normed_gauss_ds_2_update_0_stage_150 <= bright_weights_normed_gauss_ds_2_update_0_stage_149;
      bright_weights_normed_gauss_ds_2_update_0_stage_151 <= bright_weights_normed_gauss_ds_2_update_0_stage_150;
      bright_weights_normed_gauss_ds_2_update_0_stage_152 <= bright_weights_normed_gauss_ds_2_update_0_stage_151;
      bright_weights_normed_gauss_ds_2_update_0_stage_153 <= bright_weights_normed_gauss_ds_2_update_0_stage_152;
      bright_weights_normed_gauss_ds_2_update_0_stage_154 <= bright_weights_normed_gauss_ds_2_update_0_stage_153;
      bright_weights_normed_gauss_ds_2_update_0_stage_155 <= bright_weights_normed_gauss_ds_2_update_0_stage_154;
      bright_weights_normed_gauss_ds_2_update_0_stage_156 <= bright_weights_normed_gauss_ds_2_update_0_stage_155;
      bright_weights_normed_gauss_ds_2_update_0_stage_157 <= bright_weights_normed_gauss_ds_2_update_0_stage_156;
      bright_weights_normed_gauss_ds_2_update_0_stage_158 <= bright_weights_normed_gauss_ds_2_update_0_stage_157;
      bright_weights_normed_gauss_ds_2_update_0_stage_159 <= bright_weights_normed_gauss_ds_2_update_0_stage_158;
      bright_weights_normed_gauss_ds_2_update_0_stage_160 <= bright_weights_normed_gauss_ds_2_update_0_stage_159;
      bright_weights_normed_gauss_ds_2_update_0_stage_161 <= bright_weights_normed_gauss_ds_2_update_0_stage_160;
      bright_weights_normed_gauss_ds_2_update_0_stage_162 <= bright_weights_normed_gauss_ds_2_update_0_stage_161;
      bright_weights_normed_gauss_ds_2_update_0_stage_163 <= bright_weights_normed_gauss_ds_2_update_0_stage_162;
      bright_weights_normed_gauss_ds_2_update_0_stage_164 <= bright_weights_normed_gauss_ds_2_update_0_stage_163;
      bright_weights_normed_gauss_ds_2_update_0_stage_165 <= bright_weights_normed_gauss_ds_2_update_0_stage_164;
      bright_weights_normed_gauss_ds_2_update_0_stage_166 <= bright_weights_normed_gauss_ds_2_update_0_stage_165;
      bright_weights_normed_gauss_ds_2_update_0_stage_167 <= bright_weights_normed_gauss_ds_2_update_0_stage_166;
      bright_weights_normed_gauss_ds_2_update_0_stage_168 <= bright_weights_normed_gauss_ds_2_update_0_stage_167;
      bright_weights_normed_gauss_ds_2_update_0_stage_169 <= bright_weights_normed_gauss_ds_2_update_0_stage_168;
      bright_weights_normed_gauss_ds_2_update_0_stage_170 <= bright_weights_normed_gauss_ds_2_update_0_stage_169;
      bright_weights_normed_gauss_ds_2_update_0_stage_171 <= bright_weights_normed_gauss_ds_2_update_0_stage_170;
      bright_weights_normed_gauss_ds_2_update_0_stage_172 <= bright_weights_normed_gauss_ds_2_update_0_stage_171;
      bright_weights_normed_gauss_ds_2_update_0_stage_173 <= bright_weights_normed_gauss_ds_2_update_0_stage_172;
      bright_weights_normed_gauss_ds_2_update_0_stage_174 <= bright_weights_normed_gauss_ds_2_update_0_stage_173;
      bright_weights_normed_gauss_ds_2_update_0_stage_175 <= bright_weights_normed_gauss_ds_2_update_0_stage_174;
      bright_weights_normed_gauss_ds_2_update_0_stage_176 <= bright_weights_normed_gauss_ds_2_update_0_stage_175;
      bright_weights_normed_gauss_ds_2_update_0_stage_177 <= bright_weights_normed_gauss_ds_2_update_0_stage_176;
      bright_weights_normed_gauss_ds_2_update_0_stage_178 <= bright_weights_normed_gauss_ds_2_update_0_stage_177;
      bright_weights_normed_gauss_ds_2_update_0_stage_179 <= bright_weights_normed_gauss_ds_2_update_0_stage_178;
      bright_weights_normed_gauss_ds_2_update_0_stage_180 <= bright_weights_normed_gauss_ds_2_update_0_stage_179;
      bright_weights_normed_gauss_ds_2_update_0_stage_181 <= bright_weights_normed_gauss_ds_2_update_0_stage_180;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_141 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_142 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_141;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_143 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_142;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_144 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_143;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_145 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_144;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_146 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_145;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_147 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_146;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_148 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_147;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_149 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_148;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_150 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_149;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_151 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_150;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_152 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_151;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_153 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_152;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_154 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_153;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_155 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_154;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_156 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_155;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_157 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_156;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_158 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_157;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_159 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_158;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_160 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_159;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_161 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_160;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_162 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_161;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_163 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_162;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_164 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_163;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_165 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_164;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_166 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_165;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_167 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_166;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_168 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_167;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_169 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_168;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_170 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_169;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_171 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_170;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_172 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_171;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_173 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_172;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_174 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_173;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_175 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_174;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_176 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_175;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_177 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_176;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_178 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_177;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_179 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_178;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_180 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_179;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_181 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97_stage_180;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_145 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_146 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_145;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_147 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_146;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_148 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_147;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_149 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_148;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_150 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_149;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_151 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_150;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_152 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_151;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_153 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_152;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_154 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_153;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_155 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_154;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_156 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_155;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_157 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_156;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_158 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_157;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_159 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_158;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_160 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_159;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_161 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_160;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_162 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_161;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_163 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_162;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_164 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_163;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_165 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_164;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_166 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_165;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_167 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_166;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_168 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_167;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_169 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_168;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_170 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_169;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_171 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_170;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_172 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_171;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_173 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_172;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_174 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_173;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_175 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_174;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_176 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_175;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_177 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_176;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_178 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_177;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_179 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_178;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_180 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_179;
      dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_181 <= dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100_stage_180;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_146 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_147 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_146;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_148 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_147;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_149 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_148;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_150 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_149;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_151 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_150;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_152 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_151;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_153 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_152;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_154 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_153;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_155 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_154;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_156 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_155;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_157 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_156;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_158 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_157;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_159 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_158;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_160 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_159;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_161 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_160;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_162 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_161;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_163 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_162;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_164 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_163;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_165 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_164;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_166 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_165;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_167 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_166;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_168 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_167;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_169 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_168;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_170 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_169;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_171 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_170;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_172 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_171;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_173 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_172;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_174 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_173;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_175 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_174;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_176 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_175;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_177 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_176;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_178 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_177;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_179 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_178;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_180 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_179;
      dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_181 <= dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101_stage_180;
      dark_laplace_diff_2_update_0_stage_147 <= dark_laplace_diff_2_update_0;
      dark_laplace_diff_2_update_0_stage_148 <= dark_laplace_diff_2_update_0_stage_147;
      dark_laplace_diff_2_update_0_stage_149 <= dark_laplace_diff_2_update_0_stage_148;
      dark_laplace_diff_2_update_0_stage_150 <= dark_laplace_diff_2_update_0_stage_149;
      dark_laplace_diff_2_update_0_stage_151 <= dark_laplace_diff_2_update_0_stage_150;
      dark_laplace_diff_2_update_0_stage_152 <= dark_laplace_diff_2_update_0_stage_151;
      dark_laplace_diff_2_update_0_stage_153 <= dark_laplace_diff_2_update_0_stage_152;
      dark_laplace_diff_2_update_0_stage_154 <= dark_laplace_diff_2_update_0_stage_153;
      dark_laplace_diff_2_update_0_stage_155 <= dark_laplace_diff_2_update_0_stage_154;
      dark_laplace_diff_2_update_0_stage_156 <= dark_laplace_diff_2_update_0_stage_155;
      dark_laplace_diff_2_update_0_stage_157 <= dark_laplace_diff_2_update_0_stage_156;
      dark_laplace_diff_2_update_0_stage_158 <= dark_laplace_diff_2_update_0_stage_157;
      dark_laplace_diff_2_update_0_stage_159 <= dark_laplace_diff_2_update_0_stage_158;
      dark_laplace_diff_2_update_0_stage_160 <= dark_laplace_diff_2_update_0_stage_159;
      dark_laplace_diff_2_update_0_stage_161 <= dark_laplace_diff_2_update_0_stage_160;
      dark_laplace_diff_2_update_0_stage_162 <= dark_laplace_diff_2_update_0_stage_161;
      dark_laplace_diff_2_update_0_stage_163 <= dark_laplace_diff_2_update_0_stage_162;
      dark_laplace_diff_2_update_0_stage_164 <= dark_laplace_diff_2_update_0_stage_163;
      dark_laplace_diff_2_update_0_stage_165 <= dark_laplace_diff_2_update_0_stage_164;
      dark_laplace_diff_2_update_0_stage_166 <= dark_laplace_diff_2_update_0_stage_165;
      dark_laplace_diff_2_update_0_stage_167 <= dark_laplace_diff_2_update_0_stage_166;
      dark_laplace_diff_2_update_0_stage_168 <= dark_laplace_diff_2_update_0_stage_167;
      dark_laplace_diff_2_update_0_stage_169 <= dark_laplace_diff_2_update_0_stage_168;
      dark_laplace_diff_2_update_0_stage_170 <= dark_laplace_diff_2_update_0_stage_169;
      dark_laplace_diff_2_update_0_stage_171 <= dark_laplace_diff_2_update_0_stage_170;
      dark_laplace_diff_2_update_0_stage_172 <= dark_laplace_diff_2_update_0_stage_171;
      dark_laplace_diff_2_update_0_stage_173 <= dark_laplace_diff_2_update_0_stage_172;
      dark_laplace_diff_2_update_0_stage_174 <= dark_laplace_diff_2_update_0_stage_173;
      dark_laplace_diff_2_update_0_stage_175 <= dark_laplace_diff_2_update_0_stage_174;
      dark_laplace_diff_2_update_0_stage_176 <= dark_laplace_diff_2_update_0_stage_175;
      dark_laplace_diff_2_update_0_stage_177 <= dark_laplace_diff_2_update_0_stage_176;
      dark_laplace_diff_2_update_0_stage_178 <= dark_laplace_diff_2_update_0_stage_177;
      dark_laplace_diff_2_update_0_stage_179 <= dark_laplace_diff_2_update_0_stage_178;
      dark_laplace_diff_2_update_0_stage_180 <= dark_laplace_diff_2_update_0_stage_179;
      dark_laplace_diff_2_update_0_stage_181 <= dark_laplace_diff_2_update_0_stage_180;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_149 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_150 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_149;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_151 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_150;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_152 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_151;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_153 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_152;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_154 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_153;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_155 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_154;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_156 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_155;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_157 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_156;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_158 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_157;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_159 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_158;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_160 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_159;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_161 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_160;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_162 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_161;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_163 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_162;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_164 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_163;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_165 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_164;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_166 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_165;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_167 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_166;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_168 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_167;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_169 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_168;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_170 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_169;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_171 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_170;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_172 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_171;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_173 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_172;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_174 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_173;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_175 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_174;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_176 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_175;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_177 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_176;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_178 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_177;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_179 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_178;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_180 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_179;
      bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_181 <= bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103_stage_180;
      bright_weights_normed_gauss_blur_3_update_0_stage_150 <= bright_weights_normed_gauss_blur_3_update_0;
      bright_weights_normed_gauss_blur_3_update_0_stage_151 <= bright_weights_normed_gauss_blur_3_update_0_stage_150;
      bright_weights_normed_gauss_blur_3_update_0_stage_152 <= bright_weights_normed_gauss_blur_3_update_0_stage_151;
      bright_weights_normed_gauss_blur_3_update_0_stage_153 <= bright_weights_normed_gauss_blur_3_update_0_stage_152;
      bright_weights_normed_gauss_blur_3_update_0_stage_154 <= bright_weights_normed_gauss_blur_3_update_0_stage_153;
      bright_weights_normed_gauss_blur_3_update_0_stage_155 <= bright_weights_normed_gauss_blur_3_update_0_stage_154;
      bright_weights_normed_gauss_blur_3_update_0_stage_156 <= bright_weights_normed_gauss_blur_3_update_0_stage_155;
      bright_weights_normed_gauss_blur_3_update_0_stage_157 <= bright_weights_normed_gauss_blur_3_update_0_stage_156;
      bright_weights_normed_gauss_blur_3_update_0_stage_158 <= bright_weights_normed_gauss_blur_3_update_0_stage_157;
      bright_weights_normed_gauss_blur_3_update_0_stage_159 <= bright_weights_normed_gauss_blur_3_update_0_stage_158;
      bright_weights_normed_gauss_blur_3_update_0_stage_160 <= bright_weights_normed_gauss_blur_3_update_0_stage_159;
      bright_weights_normed_gauss_blur_3_update_0_stage_161 <= bright_weights_normed_gauss_blur_3_update_0_stage_160;
      bright_weights_normed_gauss_blur_3_update_0_stage_162 <= bright_weights_normed_gauss_blur_3_update_0_stage_161;
      bright_weights_normed_gauss_blur_3_update_0_stage_163 <= bright_weights_normed_gauss_blur_3_update_0_stage_162;
      bright_weights_normed_gauss_blur_3_update_0_stage_164 <= bright_weights_normed_gauss_blur_3_update_0_stage_163;
      bright_weights_normed_gauss_blur_3_update_0_stage_165 <= bright_weights_normed_gauss_blur_3_update_0_stage_164;
      bright_weights_normed_gauss_blur_3_update_0_stage_166 <= bright_weights_normed_gauss_blur_3_update_0_stage_165;
      bright_weights_normed_gauss_blur_3_update_0_stage_167 <= bright_weights_normed_gauss_blur_3_update_0_stage_166;
      bright_weights_normed_gauss_blur_3_update_0_stage_168 <= bright_weights_normed_gauss_blur_3_update_0_stage_167;
      bright_weights_normed_gauss_blur_3_update_0_stage_169 <= bright_weights_normed_gauss_blur_3_update_0_stage_168;
      bright_weights_normed_gauss_blur_3_update_0_stage_170 <= bright_weights_normed_gauss_blur_3_update_0_stage_169;
      bright_weights_normed_gauss_blur_3_update_0_stage_171 <= bright_weights_normed_gauss_blur_3_update_0_stage_170;
      bright_weights_normed_gauss_blur_3_update_0_stage_172 <= bright_weights_normed_gauss_blur_3_update_0_stage_171;
      bright_weights_normed_gauss_blur_3_update_0_stage_173 <= bright_weights_normed_gauss_blur_3_update_0_stage_172;
      bright_weights_normed_gauss_blur_3_update_0_stage_174 <= bright_weights_normed_gauss_blur_3_update_0_stage_173;
      bright_weights_normed_gauss_blur_3_update_0_stage_175 <= bright_weights_normed_gauss_blur_3_update_0_stage_174;
      bright_weights_normed_gauss_blur_3_update_0_stage_176 <= bright_weights_normed_gauss_blur_3_update_0_stage_175;
      bright_weights_normed_gauss_blur_3_update_0_stage_177 <= bright_weights_normed_gauss_blur_3_update_0_stage_176;
      bright_weights_normed_gauss_blur_3_update_0_stage_178 <= bright_weights_normed_gauss_blur_3_update_0_stage_177;
      bright_weights_normed_gauss_blur_3_update_0_stage_179 <= bright_weights_normed_gauss_blur_3_update_0_stage_178;
      bright_weights_normed_gauss_blur_3_update_0_stage_180 <= bright_weights_normed_gauss_blur_3_update_0_stage_179;
      bright_weights_normed_gauss_blur_3_update_0_stage_181 <= bright_weights_normed_gauss_blur_3_update_0_stage_180;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_151 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_152 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_151;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_153 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_152;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_154 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_153;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_155 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_154;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_156 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_155;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_157 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_156;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_158 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_157;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_159 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_158;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_160 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_159;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_161 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_160;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_162 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_161;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_163 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_162;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_164 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_163;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_165 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_164;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_166 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_165;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_167 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_166;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_168 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_167;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_169 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_168;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_170 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_169;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_171 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_170;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_172 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_171;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_173 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_172;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_174 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_173;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_175 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_174;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_176 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_175;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_177 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_176;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_178 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_177;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_179 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_178;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_180 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_179;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_181 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104_stage_180;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_152 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_153 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_152;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_154 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_153;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_155 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_154;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_156 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_155;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_157 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_156;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_158 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_157;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_159 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_158;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_160 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_159;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_161 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_160;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_162 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_161;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_163 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_162;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_164 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_163;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_165 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_164;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_166 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_165;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_167 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_166;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_168 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_167;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_169 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_168;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_170 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_169;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_171 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_170;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_172 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_171;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_173 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_172;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_174 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_173;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_175 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_174;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_176 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_175;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_177 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_176;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_178 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_177;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_179 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_178;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_180 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_179;
      bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_181 <= bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105_stage_180;
      bright_weights_normed_gauss_ds_3_update_0_stage_153 <= bright_weights_normed_gauss_ds_3_update_0;
      bright_weights_normed_gauss_ds_3_update_0_stage_154 <= bright_weights_normed_gauss_ds_3_update_0_stage_153;
      bright_weights_normed_gauss_ds_3_update_0_stage_155 <= bright_weights_normed_gauss_ds_3_update_0_stage_154;
      bright_weights_normed_gauss_ds_3_update_0_stage_156 <= bright_weights_normed_gauss_ds_3_update_0_stage_155;
      bright_weights_normed_gauss_ds_3_update_0_stage_157 <= bright_weights_normed_gauss_ds_3_update_0_stage_156;
      bright_weights_normed_gauss_ds_3_update_0_stage_158 <= bright_weights_normed_gauss_ds_3_update_0_stage_157;
      bright_weights_normed_gauss_ds_3_update_0_stage_159 <= bright_weights_normed_gauss_ds_3_update_0_stage_158;
      bright_weights_normed_gauss_ds_3_update_0_stage_160 <= bright_weights_normed_gauss_ds_3_update_0_stage_159;
      bright_weights_normed_gauss_ds_3_update_0_stage_161 <= bright_weights_normed_gauss_ds_3_update_0_stage_160;
      bright_weights_normed_gauss_ds_3_update_0_stage_162 <= bright_weights_normed_gauss_ds_3_update_0_stage_161;
      bright_weights_normed_gauss_ds_3_update_0_stage_163 <= bright_weights_normed_gauss_ds_3_update_0_stage_162;
      bright_weights_normed_gauss_ds_3_update_0_stage_164 <= bright_weights_normed_gauss_ds_3_update_0_stage_163;
      bright_weights_normed_gauss_ds_3_update_0_stage_165 <= bright_weights_normed_gauss_ds_3_update_0_stage_164;
      bright_weights_normed_gauss_ds_3_update_0_stage_166 <= bright_weights_normed_gauss_ds_3_update_0_stage_165;
      bright_weights_normed_gauss_ds_3_update_0_stage_167 <= bright_weights_normed_gauss_ds_3_update_0_stage_166;
      bright_weights_normed_gauss_ds_3_update_0_stage_168 <= bright_weights_normed_gauss_ds_3_update_0_stage_167;
      bright_weights_normed_gauss_ds_3_update_0_stage_169 <= bright_weights_normed_gauss_ds_3_update_0_stage_168;
      bright_weights_normed_gauss_ds_3_update_0_stage_170 <= bright_weights_normed_gauss_ds_3_update_0_stage_169;
      bright_weights_normed_gauss_ds_3_update_0_stage_171 <= bright_weights_normed_gauss_ds_3_update_0_stage_170;
      bright_weights_normed_gauss_ds_3_update_0_stage_172 <= bright_weights_normed_gauss_ds_3_update_0_stage_171;
      bright_weights_normed_gauss_ds_3_update_0_stage_173 <= bright_weights_normed_gauss_ds_3_update_0_stage_172;
      bright_weights_normed_gauss_ds_3_update_0_stage_174 <= bright_weights_normed_gauss_ds_3_update_0_stage_173;
      bright_weights_normed_gauss_ds_3_update_0_stage_175 <= bright_weights_normed_gauss_ds_3_update_0_stage_174;
      bright_weights_normed_gauss_ds_3_update_0_stage_176 <= bright_weights_normed_gauss_ds_3_update_0_stage_175;
      bright_weights_normed_gauss_ds_3_update_0_stage_177 <= bright_weights_normed_gauss_ds_3_update_0_stage_176;
      bright_weights_normed_gauss_ds_3_update_0_stage_178 <= bright_weights_normed_gauss_ds_3_update_0_stage_177;
      bright_weights_normed_gauss_ds_3_update_0_stage_179 <= bright_weights_normed_gauss_ds_3_update_0_stage_178;
      bright_weights_normed_gauss_ds_3_update_0_stage_180 <= bright_weights_normed_gauss_ds_3_update_0_stage_179;
      bright_weights_normed_gauss_ds_3_update_0_stage_181 <= bright_weights_normed_gauss_ds_3_update_0_stage_180;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_155 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_156 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_155;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_157 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_156;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_158 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_157;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_159 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_158;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_160 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_159;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_161 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_160;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_162 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_161;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_163 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_162;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_164 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_163;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_165 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_164;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_166 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_165;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_167 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_166;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_168 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_167;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_169 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_168;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_170 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_169;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_171 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_170;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_172 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_171;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_173 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_172;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_174 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_173;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_175 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_174;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_176 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_175;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_177 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_176;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_178 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_177;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_179 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_178;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_180 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_179;
      bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_181 <= bright_laplace_diff_2_fused_level_2_update_0_read_read_107_stage_180;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_154 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_155 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_154;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_156 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_155;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_157 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_156;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_158 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_157;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_159 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_158;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_160 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_159;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_161 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_160;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_162 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_161;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_163 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_162;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_164 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_163;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_165 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_164;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_166 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_165;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_167 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_166;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_168 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_167;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_169 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_168;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_170 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_169;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_171 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_170;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_172 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_171;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_173 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_172;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_174 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_173;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_175 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_174;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_176 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_175;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_177 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_176;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_178 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_177;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_179 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_178;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_180 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_179;
      bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_181 <= bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106_stage_180;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_156 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_157 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_156;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_158 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_157;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_159 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_158;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_160 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_159;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_161 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_160;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_162 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_161;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_163 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_162;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_164 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_163;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_165 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_164;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_166 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_165;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_167 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_166;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_168 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_167;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_169 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_168;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_170 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_169;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_171 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_170;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_172 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_171;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_173 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_172;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_174 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_173;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_175 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_174;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_176 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_175;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_177 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_176;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_178 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_177;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_179 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_178;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_180 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_179;
      dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_181 <= dark_laplace_diff_2_fused_level_2_update_0_read_read_108_stage_180;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_157 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_158 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_157;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_159 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_158;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_160 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_159;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_161 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_160;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_162 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_161;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_163 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_162;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_164 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_163;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_165 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_164;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_166 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_165;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_167 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_166;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_168 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_167;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_169 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_168;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_170 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_169;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_171 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_170;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_172 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_171;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_173 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_172;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_174 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_173;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_175 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_174;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_176 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_175;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_177 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_176;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_178 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_177;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_179 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_178;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_180 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_179;
      bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_181 <= bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109_stage_180;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_158 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_159 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_158;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_160 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_159;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_161 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_160;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_162 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_161;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_163 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_162;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_164 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_163;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_165 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_164;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_166 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_165;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_167 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_166;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_168 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_167;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_169 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_168;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_170 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_169;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_171 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_170;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_172 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_171;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_173 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_172;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_174 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_173;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_175 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_174;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_176 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_175;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_177 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_176;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_178 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_177;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_179 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_178;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_180 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_179;
      dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_181 <= dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110_stage_180;
      fused_level_2_update_0_stage_159 <= fused_level_2_update_0;
      fused_level_2_update_0_stage_160 <= fused_level_2_update_0_stage_159;
      fused_level_2_update_0_stage_161 <= fused_level_2_update_0_stage_160;
      fused_level_2_update_0_stage_162 <= fused_level_2_update_0_stage_161;
      fused_level_2_update_0_stage_163 <= fused_level_2_update_0_stage_162;
      fused_level_2_update_0_stage_164 <= fused_level_2_update_0_stage_163;
      fused_level_2_update_0_stage_165 <= fused_level_2_update_0_stage_164;
      fused_level_2_update_0_stage_166 <= fused_level_2_update_0_stage_165;
      fused_level_2_update_0_stage_167 <= fused_level_2_update_0_stage_166;
      fused_level_2_update_0_stage_168 <= fused_level_2_update_0_stage_167;
      fused_level_2_update_0_stage_169 <= fused_level_2_update_0_stage_168;
      fused_level_2_update_0_stage_170 <= fused_level_2_update_0_stage_169;
      fused_level_2_update_0_stage_171 <= fused_level_2_update_0_stage_170;
      fused_level_2_update_0_stage_172 <= fused_level_2_update_0_stage_171;
      fused_level_2_update_0_stage_173 <= fused_level_2_update_0_stage_172;
      fused_level_2_update_0_stage_174 <= fused_level_2_update_0_stage_173;
      fused_level_2_update_0_stage_175 <= fused_level_2_update_0_stage_174;
      fused_level_2_update_0_stage_176 <= fused_level_2_update_0_stage_175;
      fused_level_2_update_0_stage_177 <= fused_level_2_update_0_stage_176;
      fused_level_2_update_0_stage_178 <= fused_level_2_update_0_stage_177;
      fused_level_2_update_0_stage_179 <= fused_level_2_update_0_stage_178;
      fused_level_2_update_0_stage_180 <= fused_level_2_update_0_stage_179;
      fused_level_2_update_0_stage_181 <= fused_level_2_update_0_stage_180;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_160 <= fused_level_2_fused_level_2_update_0_write_write_111;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_161 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_160;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_162 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_161;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_163 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_162;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_164 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_163;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_165 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_164;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_166 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_165;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_167 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_166;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_168 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_167;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_169 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_168;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_170 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_169;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_171 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_170;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_172 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_171;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_173 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_172;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_174 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_173;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_175 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_174;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_176 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_175;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_177 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_176;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_178 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_177;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_179 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_178;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_180 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_179;
      fused_level_2_fused_level_2_update_0_write_write_111_stage_181 <= fused_level_2_fused_level_2_update_0_write_write_111_stage_180;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_161 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_162 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_161;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_163 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_162;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_164 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_163;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_165 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_164;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_166 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_165;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_167 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_166;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_168 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_167;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_169 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_168;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_170 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_169;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_171 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_170;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_172 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_171;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_173 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_172;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_174 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_173;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_175 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_174;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_176 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_175;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_177 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_176;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_178 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_177;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_179 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_178;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_180 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_179;
      bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_181 <= bright_gauss_ds_3_fused_level_3_update_0_read_read_112_stage_180;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_162 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_163 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_162;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_164 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_163;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_165 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_164;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_166 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_165;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_167 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_166;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_168 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_167;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_169 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_168;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_170 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_169;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_171 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_170;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_172 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_171;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_173 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_172;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_174 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_173;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_175 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_174;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_176 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_175;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_177 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_176;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_178 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_177;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_179 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_178;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_180 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_179;
      dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_181 <= dark_gauss_ds_3_fused_level_3_update_0_read_read_113_stage_180;


    end

  end


  // Data processing units...
  // buf_bright_gauss_blur_1
  logic [0:0] buf_bright_gauss_blur_1_clk;
  logic [0:0] buf_bright_gauss_blur_1_rst;
  logic [0:0] buf_bright_gauss_blur_1_start;
  logic [0:0] buf_bright_gauss_blur_1_done;
  logic [0:0] buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wen;
  logic [31:0] buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wdata;
  logic [31:0] buf_bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_rdata;
  bright_gauss_blur_1 buf_bright_gauss_blur_1(.clk(buf_bright_gauss_blur_1_clk), .rst(buf_bright_gauss_blur_1_rst), .start(buf_bright_gauss_blur_1_start), .done(buf_bright_gauss_blur_1_done), .bright_gauss_blur_1_update_0_write_wen(buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wen), .bright_gauss_blur_1_update_0_write_wdata(buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wdata), .bright_gauss_ds_1_update_0_read_dummy(buf_bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_dummy), .bright_gauss_ds_1_update_0_read_rdata(buf_bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_rdata));
  assign buf_bright_gauss_blur_1_clk = clk;
  assign buf_bright_gauss_blur_1_rst = rst;
  assign buf_bright_gauss_blur_1_start = start;
  // Bindings to buf_bright_gauss_blur_1
    // bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13
  assign bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_write_13 = buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wdata;
  assign buf_bright_gauss_blur_1_bright_gauss_blur_1_update_0_write_wen = stage_20_active;
    // bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20
  assign bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_read_20 = buf_bright_gauss_blur_1_bright_gauss_ds_1_update_0_read_rdata;

  // buf_bright_gauss_blur_2
  logic [0:0] buf_bright_gauss_blur_2_clk;
  logic [0:0] buf_bright_gauss_blur_2_rst;
  logic [0:0] buf_bright_gauss_blur_2_start;
  logic [0:0] buf_bright_gauss_blur_2_done;
  logic [0:0] buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wen;
  logic [31:0] buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wdata;
  logic [31:0] buf_bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_rdata;
  bright_gauss_blur_2 buf_bright_gauss_blur_2(.clk(buf_bright_gauss_blur_2_clk), .rst(buf_bright_gauss_blur_2_rst), .start(buf_bright_gauss_blur_2_start), .done(buf_bright_gauss_blur_2_done), .bright_gauss_blur_2_update_0_write_wen(buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wen), .bright_gauss_blur_2_update_0_write_wdata(buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wdata), .bright_gauss_ds_2_update_0_read_dummy(buf_bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_dummy), .bright_gauss_ds_2_update_0_read_rdata(buf_bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_rdata));
  assign buf_bright_gauss_blur_2_clk = clk;
  assign buf_bright_gauss_blur_2_rst = rst;
  assign buf_bright_gauss_blur_2_start = start;
  // Bindings to buf_bright_gauss_blur_2
    // bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32
  assign bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_read_32 = buf_bright_gauss_blur_2_bright_gauss_ds_2_update_0_read_rdata;
    // bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26
  assign bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_write_26 = buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wdata;
  assign buf_bright_gauss_blur_2_bright_gauss_blur_2_update_0_write_wen = stage_39_active;

  // buf_bright
  logic [0:0] buf_bright_clk;
  logic [0:0] buf_bright_rst;
  logic [0:0] buf_bright_start;
  logic [0:0] buf_bright_done;
  logic [0:0] buf_bright_bright_update_0_write_wen;
  logic [31:0] buf_bright_bright_weights_update_0_read_dummy;
  logic [31:0] buf_bright_bright_update_0_write_wdata;
  logic [287:0] buf_bright_bright_gauss_blur_1_update_0_read_dummy;
  logic [287:0] buf_bright_bright_gauss_blur_1_update_0_read_rdata;
  logic [31:0] buf_bright_bright_laplace_diff_0_update_0_read_dummy;
  logic [31:0] buf_bright_bright_laplace_diff_0_update_0_read_rdata;
  logic [31:0] buf_bright_bright_weights_update_0_read_rdata;
  bright buf_bright(.clk(buf_bright_clk), .rst(buf_bright_rst), .start(buf_bright_start), .done(buf_bright_done), .bright_update_0_write_wen(buf_bright_bright_update_0_write_wen), .bright_weights_update_0_read_dummy(buf_bright_bright_weights_update_0_read_dummy), .bright_update_0_write_wdata(buf_bright_bright_update_0_write_wdata), .bright_gauss_blur_1_update_0_read_dummy(buf_bright_bright_gauss_blur_1_update_0_read_dummy), .bright_gauss_blur_1_update_0_read_rdata(buf_bright_bright_gauss_blur_1_update_0_read_rdata), .bright_laplace_diff_0_update_0_read_dummy(buf_bright_bright_laplace_diff_0_update_0_read_dummy), .bright_laplace_diff_0_update_0_read_rdata(buf_bright_bright_laplace_diff_0_update_0_read_rdata), .bright_weights_update_0_read_rdata(buf_bright_bright_weights_update_0_read_rdata));
  assign buf_bright_clk = clk;
  assign buf_bright_rst = rst;
  assign buf_bright_start = start;
  // Bindings to buf_bright
    // bright_bright_weights_update_0_read_read_4
  assign bright_bright_weights_update_0_read_read_4 = buf_bright_bright_weights_update_0_read_rdata;
    // bright_bright_update_0_write_write_3
  assign bright_bright_update_0_write_write_3 = buf_bright_bright_update_0_write_wdata;
  assign buf_bright_bright_update_0_write_wen = stage_5_active;
    // bright_bright_gauss_blur_1_update_0_read_read_12
  assign bright_bright_gauss_blur_1_update_0_read_read_12 = buf_bright_bright_gauss_blur_1_update_0_read_rdata;
    // bright_bright_laplace_diff_0_update_0_read_read_42
  assign bright_bright_laplace_diff_0_update_0_read_read_42 = buf_bright_bright_laplace_diff_0_update_0_read_rdata;

  // buf_bright_gauss_ds_1
  logic [0:0] buf_bright_gauss_ds_1_clk;
  logic [0:0] buf_bright_gauss_ds_1_rst;
  logic [0:0] buf_bright_gauss_ds_1_start;
  logic [0:0] buf_bright_gauss_ds_1_done;
  logic [287:0] buf_bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_dummy;
  logic [0:0] buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wen;
  logic [31:0] buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wdata;
  logic [287:0] buf_bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_rdata;
  logic [31:0] buf_bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_rdata;
  logic [31:0] buf_bright_gauss_ds_1_bright_laplace_us_0_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_ds_1_bright_laplace_us_0_update_0_read_rdata;
  bright_gauss_ds_1 buf_bright_gauss_ds_1(.clk(buf_bright_gauss_ds_1_clk), .rst(buf_bright_gauss_ds_1_rst), .start(buf_bright_gauss_ds_1_start), .done(buf_bright_gauss_ds_1_done), .bright_gauss_blur_2_update_0_read_dummy(buf_bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_dummy), .bright_gauss_ds_1_update_0_write_wen(buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wen), .bright_gauss_ds_1_update_0_write_wdata(buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wdata), .bright_gauss_blur_2_update_0_read_rdata(buf_bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_rdata), .bright_laplace_diff_1_update_0_read_dummy(buf_bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_dummy), .bright_laplace_diff_1_update_0_read_rdata(buf_bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_rdata), .bright_laplace_us_0_update_0_read_dummy(buf_bright_gauss_ds_1_bright_laplace_us_0_update_0_read_dummy), .bright_laplace_us_0_update_0_read_rdata(buf_bright_gauss_ds_1_bright_laplace_us_0_update_0_read_rdata));
  assign buf_bright_gauss_ds_1_clk = clk;
  assign buf_bright_gauss_ds_1_rst = rst;
  assign buf_bright_gauss_ds_1_start = start;
  // Bindings to buf_bright_gauss_ds_1
    // bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21
  assign bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_write_21 = buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wdata;
  assign buf_bright_gauss_ds_1_bright_gauss_ds_1_update_0_write_wen = stage_32_active;
    // bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25
  assign bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_read_25 = buf_bright_gauss_ds_1_bright_gauss_blur_2_update_0_read_rdata;
    // bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30
  assign bright_gauss_ds_1_bright_laplace_us_0_update_0_read_read_30 = buf_bright_gauss_ds_1_bright_laplace_us_0_update_0_read_rdata;
    // bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67
  assign bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_read_67 = buf_bright_gauss_ds_1_bright_laplace_diff_1_update_0_read_rdata;

  // buf_bright_gauss_blur_3
  logic [0:0] buf_bright_gauss_blur_3_clk;
  logic [0:0] buf_bright_gauss_blur_3_rst;
  logic [0:0] buf_bright_gauss_blur_3_start;
  logic [0:0] buf_bright_gauss_blur_3_done;
  logic [0:0] buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wen;
  logic [31:0] buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wdata;
  logic [31:0] buf_bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_rdata;
  bright_gauss_blur_3 buf_bright_gauss_blur_3(.clk(buf_bright_gauss_blur_3_clk), .rst(buf_bright_gauss_blur_3_rst), .start(buf_bright_gauss_blur_3_start), .done(buf_bright_gauss_blur_3_done), .bright_gauss_blur_3_update_0_write_wen(buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wen), .bright_gauss_blur_3_update_0_write_wdata(buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wdata), .bright_gauss_ds_3_update_0_read_dummy(buf_bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_dummy), .bright_gauss_ds_3_update_0_read_rdata(buf_bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_rdata));
  assign buf_bright_gauss_blur_3_clk = clk;
  assign buf_bright_gauss_blur_3_rst = rst;
  assign buf_bright_gauss_blur_3_start = start;
  // Bindings to buf_bright_gauss_blur_3
    // bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38
  assign bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_read_38 = buf_bright_gauss_blur_3_bright_gauss_ds_3_update_0_read_rdata;
    // bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37
  assign bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_write_37 = buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wdata;
  assign buf_bright_gauss_blur_3_bright_gauss_blur_3_update_0_write_wen = stage_55_active;

  // buf_bright_gauss_ds_2
  logic [0:0] buf_bright_gauss_ds_2_clk;
  logic [0:0] buf_bright_gauss_ds_2_rst;
  logic [0:0] buf_bright_gauss_ds_2_start;
  logic [0:0] buf_bright_gauss_ds_2_done;
  logic [0:0] buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wen;
  logic [31:0] buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wdata;
  logic [287:0] buf_bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_dummy;
  logic [287:0] buf_bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_rdata;
  logic [31:0] buf_bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_rdata;
  logic [31:0] buf_bright_gauss_ds_2_bright_laplace_us_1_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_ds_2_bright_laplace_us_1_update_0_read_rdata;
  bright_gauss_ds_2 buf_bright_gauss_ds_2(.clk(buf_bright_gauss_ds_2_clk), .rst(buf_bright_gauss_ds_2_rst), .start(buf_bright_gauss_ds_2_start), .done(buf_bright_gauss_ds_2_done), .bright_gauss_ds_2_update_0_write_wen(buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wen), .bright_gauss_ds_2_update_0_write_wdata(buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wdata), .bright_gauss_blur_3_update_0_read_dummy(buf_bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_dummy), .bright_gauss_blur_3_update_0_read_rdata(buf_bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_rdata), .bright_laplace_diff_2_update_0_read_dummy(buf_bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_dummy), .bright_laplace_diff_2_update_0_read_rdata(buf_bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_rdata), .bright_laplace_us_1_update_0_read_dummy(buf_bright_gauss_ds_2_bright_laplace_us_1_update_0_read_dummy), .bright_laplace_us_1_update_0_read_rdata(buf_bright_gauss_ds_2_bright_laplace_us_1_update_0_read_rdata));
  assign buf_bright_gauss_ds_2_clk = clk;
  assign buf_bright_gauss_ds_2_rst = rst;
  assign buf_bright_gauss_ds_2_start = start;
  // Bindings to buf_bright_gauss_ds_2
    // bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40
  assign bright_gauss_ds_2_bright_laplace_us_1_update_0_read_read_40 = buf_bright_gauss_ds_2_bright_laplace_us_1_update_0_read_rdata;
    // bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33
  assign bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_write_33 = buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wdata;
  assign buf_bright_gauss_ds_2_bright_gauss_ds_2_update_0_write_wen = stage_49_active;
    // bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36
  assign bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_read_36 = buf_bright_gauss_ds_2_bright_gauss_blur_3_update_0_read_rdata;
    // bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82
  assign bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_read_82 = buf_bright_gauss_ds_2_bright_laplace_diff_2_update_0_read_rdata;

  // buf_bright_gauss_ds_3
  logic [0:0] buf_bright_gauss_ds_3_clk;
  logic [0:0] buf_bright_gauss_ds_3_rst;
  logic [0:0] buf_bright_gauss_ds_3_start;
  logic [0:0] buf_bright_gauss_ds_3_done;
  logic [31:0] buf_bright_gauss_ds_3_fused_level_3_update_0_read_dummy;
  logic [0:0] buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wen;
  logic [31:0] buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wdata;
  logic [31:0] buf_bright_gauss_ds_3_bright_laplace_us_2_update_0_read_dummy;
  logic [31:0] buf_bright_gauss_ds_3_bright_laplace_us_2_update_0_read_rdata;
  logic [31:0] buf_bright_gauss_ds_3_fused_level_3_update_0_read_rdata;
  bright_gauss_ds_3 buf_bright_gauss_ds_3(.clk(buf_bright_gauss_ds_3_clk), .rst(buf_bright_gauss_ds_3_rst), .start(buf_bright_gauss_ds_3_start), .done(buf_bright_gauss_ds_3_done), .fused_level_3_update_0_read_dummy(buf_bright_gauss_ds_3_fused_level_3_update_0_read_dummy), .bright_gauss_ds_3_update_0_write_wen(buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wen), .bright_gauss_ds_3_update_0_write_wdata(buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wdata), .bright_laplace_us_2_update_0_read_dummy(buf_bright_gauss_ds_3_bright_laplace_us_2_update_0_read_dummy), .bright_laplace_us_2_update_0_read_rdata(buf_bright_gauss_ds_3_bright_laplace_us_2_update_0_read_rdata), .fused_level_3_update_0_read_rdata(buf_bright_gauss_ds_3_fused_level_3_update_0_read_rdata));
  assign buf_bright_gauss_ds_3_clk = clk;
  assign buf_bright_gauss_ds_3_rst = rst;
  assign buf_bright_gauss_ds_3_start = start;
  // Bindings to buf_bright_gauss_ds_3
    // bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39
  assign bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_write_39 = buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wdata;
  assign buf_bright_gauss_ds_3_bright_gauss_ds_3_update_0_write_wen = stage_58_active;
    // bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59
  assign bright_gauss_ds_3_bright_laplace_us_2_update_0_read_read_59 = buf_bright_gauss_ds_3_bright_laplace_us_2_update_0_read_rdata;
    // bright_gauss_ds_3_fused_level_3_update_0_read_read_112
  assign bright_gauss_ds_3_fused_level_3_update_0_read_read_112 = buf_bright_gauss_ds_3_fused_level_3_update_0_read_rdata;

  // buf_bright_laplace_diff_0
  logic [0:0] buf_bright_laplace_diff_0_clk;
  logic [0:0] buf_bright_laplace_diff_0_rst;
  logic [0:0] buf_bright_laplace_diff_0_start;
  logic [0:0] buf_bright_laplace_diff_0_done;
  logic [0:0] buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wen;
  logic [31:0] buf_bright_laplace_diff_0_fused_level_0_update_0_read_dummy;
  logic [31:0] buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_diff_0_fused_level_0_update_0_read_rdata;
  bright_laplace_diff_0 buf_bright_laplace_diff_0(.clk(buf_bright_laplace_diff_0_clk), .rst(buf_bright_laplace_diff_0_rst), .start(buf_bright_laplace_diff_0_start), .done(buf_bright_laplace_diff_0_done), .bright_laplace_diff_0_update_0_write_wen(buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wen), .fused_level_0_update_0_read_dummy(buf_bright_laplace_diff_0_fused_level_0_update_0_read_dummy), .bright_laplace_diff_0_update_0_write_wdata(buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wdata), .fused_level_0_update_0_read_rdata(buf_bright_laplace_diff_0_fused_level_0_update_0_read_rdata));
  assign buf_bright_laplace_diff_0_clk = clk;
  assign buf_bright_laplace_diff_0_rst = rst;
  assign buf_bright_laplace_diff_0_start = start;
  // Bindings to buf_bright_laplace_diff_0
    // bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44
  assign bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_write_44 = buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wdata;
  assign buf_bright_laplace_diff_0_bright_laplace_diff_0_update_0_write_wen = stage_65_active;
    // bright_laplace_diff_0_fused_level_0_update_0_read_read_77
  assign bright_laplace_diff_0_fused_level_0_update_0_read_read_77 = buf_bright_laplace_diff_0_fused_level_0_update_0_read_rdata;

  // buf_bright_laplace_diff_1
  logic [0:0] buf_bright_laplace_diff_1_clk;
  logic [0:0] buf_bright_laplace_diff_1_rst;
  logic [0:0] buf_bright_laplace_diff_1_start;
  logic [0:0] buf_bright_laplace_diff_1_done;
  logic [31:0] buf_bright_laplace_diff_1_fused_level_1_update_0_read_dummy;
  logic [0:0] buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wen;
  logic [31:0] buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_diff_1_fused_level_1_update_0_read_rdata;
  bright_laplace_diff_1 buf_bright_laplace_diff_1(.clk(buf_bright_laplace_diff_1_clk), .rst(buf_bright_laplace_diff_1_rst), .start(buf_bright_laplace_diff_1_start), .done(buf_bright_laplace_diff_1_done), .fused_level_1_update_0_read_dummy(buf_bright_laplace_diff_1_fused_level_1_update_0_read_dummy), .bright_laplace_diff_1_update_0_write_wen(buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wen), .bright_laplace_diff_1_update_0_write_wdata(buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wdata), .fused_level_1_update_0_read_rdata(buf_bright_laplace_diff_1_fused_level_1_update_0_read_rdata));
  assign buf_bright_laplace_diff_1_clk = clk;
  assign buf_bright_laplace_diff_1_rst = rst;
  assign buf_bright_laplace_diff_1_start = start;
  // Bindings to buf_bright_laplace_diff_1
    // bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69
  assign bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_write_69 = buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wdata;
  assign buf_bright_laplace_diff_1_bright_laplace_diff_1_update_0_write_wen = stage_101_active;
    // bright_laplace_diff_1_fused_level_1_update_0_read_read_85
  assign bright_laplace_diff_1_fused_level_1_update_0_read_read_85 = buf_bright_laplace_diff_1_fused_level_1_update_0_read_rdata;

  // bright_laplace_us_1_update_0_137
  logic [0:0] bright_laplace_us_1_update_0_137_clk;
  logic [0:0] bright_laplace_us_1_update_0_137_rst;
  logic [0:0] bright_laplace_us_1_update_0_137_start;
  logic [0:0] bright_laplace_us_1_update_0_137_done;
  logic [31:0] bright_laplace_us_1_update_0_137_src_in;
  logic [31:0] bright_laplace_us_1_update_0_137_src_out;
  logic [31:0] bright_laplace_us_1_update_0_137_out;
  bright_laplace_us_1_update_0 bright_laplace_us_1_update_0_137(.clk(bright_laplace_us_1_update_0_137_clk), .rst(bright_laplace_us_1_update_0_137_rst), .start(bright_laplace_us_1_update_0_137_start), .done(bright_laplace_us_1_update_0_137_done), .src_in(bright_laplace_us_1_update_0_137_src_in), .src_out(bright_laplace_us_1_update_0_137_src_out), .out(bright_laplace_us_1_update_0_137_out));
  assign bright_laplace_us_1_update_0_137_clk = clk;
  assign bright_laplace_us_1_update_0_137_rst = rst;
  assign bright_laplace_us_1_update_0_137_start = start;
  // Bindings to bright_laplace_us_1_update_0_137
    // bright_laplace_us_1_update_0
  assign bright_laplace_us_1_update_0 = bright_laplace_us_1_update_0_137_out;

  // weight_sums_update_0_144
  logic [0:0] weight_sums_update_0_144_clk;
  logic [0:0] weight_sums_update_0_144_rst;
  logic [0:0] weight_sums_update_0_144_start;
  logic [0:0] weight_sums_update_0_144_done;
  logic [31:0] weight_sums_update_0_144_src_in;
  logic [31:0] weight_sums_update_0_144_src_out;
  logic [31:0] weight_sums_update_0_144_out;
  weight_sums_update_0 weight_sums_update_0_144(.clk(weight_sums_update_0_144_clk), .rst(weight_sums_update_0_144_rst), .start(weight_sums_update_0_144_start), .done(weight_sums_update_0_144_done), .src_in(weight_sums_update_0_144_src_in), .src_out(weight_sums_update_0_144_src_out), .out(weight_sums_update_0_144_out));
  assign weight_sums_update_0_144_clk = clk;
  assign weight_sums_update_0_144_rst = rst;
  assign weight_sums_update_0_144_start = start;
  // Bindings to weight_sums_update_0_144
    // weight_sums_update_0
  assign weight_sums_update_0 = weight_sums_update_0_144_out;

  // dark_laplace_us_0_update_0_143
  logic [0:0] dark_laplace_us_0_update_0_143_clk;
  logic [0:0] dark_laplace_us_0_update_0_143_rst;
  logic [0:0] dark_laplace_us_0_update_0_143_start;
  logic [0:0] dark_laplace_us_0_update_0_143_done;
  logic [31:0] dark_laplace_us_0_update_0_143_src_in;
  logic [31:0] dark_laplace_us_0_update_0_143_src_out;
  logic [31:0] dark_laplace_us_0_update_0_143_out;
  dark_laplace_us_0_update_0 dark_laplace_us_0_update_0_143(.clk(dark_laplace_us_0_update_0_143_clk), .rst(dark_laplace_us_0_update_0_143_rst), .start(dark_laplace_us_0_update_0_143_start), .done(dark_laplace_us_0_update_0_143_done), .src_in(dark_laplace_us_0_update_0_143_src_in), .src_out(dark_laplace_us_0_update_0_143_src_out), .out(dark_laplace_us_0_update_0_143_out));
  assign dark_laplace_us_0_update_0_143_clk = clk;
  assign dark_laplace_us_0_update_0_143_rst = rst;
  assign dark_laplace_us_0_update_0_143_start = start;
  // Bindings to dark_laplace_us_0_update_0_143
    // dark_laplace_us_0_update_0
  assign dark_laplace_us_0_update_0 = dark_laplace_us_0_update_0_143_out;

  // fused_level_3_update_0_140
  logic [0:0] fused_level_3_update_0_140_clk;
  logic [0:0] fused_level_3_update_0_140_rst;
  logic [0:0] fused_level_3_update_0_140_start;
  logic [0:0] fused_level_3_update_0_140_done;
  logic [31:0] fused_level_3_update_0_140_src_in;
  logic [31:0] fused_level_3_update_0_140_src_out;
  logic [31:0] fused_level_3_update_0_140_out;
  fused_level_3_update_0 fused_level_3_update_0_140(.clk(fused_level_3_update_0_140_clk), .rst(fused_level_3_update_0_140_rst), .start(fused_level_3_update_0_140_start), .done(fused_level_3_update_0_140_done), .src_in(fused_level_3_update_0_140_src_in), .src_out(fused_level_3_update_0_140_src_out), .out(fused_level_3_update_0_140_out));
  assign fused_level_3_update_0_140_clk = clk;
  assign fused_level_3_update_0_140_rst = rst;
  assign fused_level_3_update_0_140_start = start;
  // Bindings to fused_level_3_update_0_140
    // fused_level_3_update_0
  assign fused_level_3_update_0 = fused_level_3_update_0_140_out;

  // final_merged_0_update_0_142
  logic [0:0] final_merged_0_update_0_142_clk;
  logic [0:0] final_merged_0_update_0_142_rst;
  logic [0:0] final_merged_0_update_0_142_start;
  logic [0:0] final_merged_0_update_0_142_done;
  logic [31:0] final_merged_0_update_0_142_src_in;
  logic [31:0] final_merged_0_update_0_142_src_out;
  logic [31:0] final_merged_0_update_0_142_out;
  final_merged_0_update_0 final_merged_0_update_0_142(.clk(final_merged_0_update_0_142_clk), .rst(final_merged_0_update_0_142_rst), .start(final_merged_0_update_0_142_start), .done(final_merged_0_update_0_142_done), .src_in(final_merged_0_update_0_142_src_in), .src_out(final_merged_0_update_0_142_src_out), .out(final_merged_0_update_0_142_out));
  assign final_merged_0_update_0_142_clk = clk;
  assign final_merged_0_update_0_142_rst = rst;
  assign final_merged_0_update_0_142_start = start;
  // Bindings to final_merged_0_update_0_142
    // final_merged_0_update_0
  assign final_merged_0_update_0 = final_merged_0_update_0_142_out;

  // dark_laplace_diff_0_update_0_145
  logic [0:0] dark_laplace_diff_0_update_0_145_clk;
  logic [0:0] dark_laplace_diff_0_update_0_145_rst;
  logic [0:0] dark_laplace_diff_0_update_0_145_start;
  logic [0:0] dark_laplace_diff_0_update_0_145_done;
  logic [31:0] dark_laplace_diff_0_update_0_145_src_in;
  logic [31:0] dark_laplace_diff_0_update_0_145_src_out;
  logic [31:0] dark_laplace_diff_0_update_0_145_out;
  dark_laplace_diff_0_update_0 dark_laplace_diff_0_update_0_145(.clk(dark_laplace_diff_0_update_0_145_clk), .rst(dark_laplace_diff_0_update_0_145_rst), .start(dark_laplace_diff_0_update_0_145_start), .done(dark_laplace_diff_0_update_0_145_done), .src_in(dark_laplace_diff_0_update_0_145_src_in), .src_out(dark_laplace_diff_0_update_0_145_src_out), .out(dark_laplace_diff_0_update_0_145_out));
  assign dark_laplace_diff_0_update_0_145_clk = clk;
  assign dark_laplace_diff_0_update_0_145_rst = rst;
  assign dark_laplace_diff_0_update_0_145_start = start;
  // Bindings to dark_laplace_diff_0_update_0_145
    // dark_laplace_diff_0_update_0
  assign dark_laplace_diff_0_update_0 = dark_laplace_diff_0_update_0_145_out;

  // bright_laplace_us_2_update_0_139
  logic [0:0] bright_laplace_us_2_update_0_139_clk;
  logic [0:0] bright_laplace_us_2_update_0_139_rst;
  logic [0:0] bright_laplace_us_2_update_0_139_start;
  logic [0:0] bright_laplace_us_2_update_0_139_done;
  logic [31:0] bright_laplace_us_2_update_0_139_src_in;
  logic [31:0] bright_laplace_us_2_update_0_139_src_out;
  logic [31:0] bright_laplace_us_2_update_0_139_out;
  bright_laplace_us_2_update_0 bright_laplace_us_2_update_0_139(.clk(bright_laplace_us_2_update_0_139_clk), .rst(bright_laplace_us_2_update_0_139_rst), .start(bright_laplace_us_2_update_0_139_start), .done(bright_laplace_us_2_update_0_139_done), .src_in(bright_laplace_us_2_update_0_139_src_in), .src_out(bright_laplace_us_2_update_0_139_src_out), .out(bright_laplace_us_2_update_0_139_out));
  assign bright_laplace_us_2_update_0_139_clk = clk;
  assign bright_laplace_us_2_update_0_139_rst = rst;
  assign bright_laplace_us_2_update_0_139_start = start;
  // Bindings to bright_laplace_us_2_update_0_139
    // bright_laplace_us_2_update_0
  assign bright_laplace_us_2_update_0 = bright_laplace_us_2_update_0_139_out;

  // dark_weights_normed_gauss_ds_1_update_0_150
  logic [0:0] dark_weights_normed_gauss_ds_1_update_0_150_clk;
  logic [0:0] dark_weights_normed_gauss_ds_1_update_0_150_rst;
  logic [0:0] dark_weights_normed_gauss_ds_1_update_0_150_start;
  logic [0:0] dark_weights_normed_gauss_ds_1_update_0_150_done;
  logic [31:0] dark_weights_normed_gauss_ds_1_update_0_150_src_in;
  logic [31:0] dark_weights_normed_gauss_ds_1_update_0_150_src_out;
  logic [31:0] dark_weights_normed_gauss_ds_1_update_0_150_out;
  dark_weights_normed_gauss_ds_1_update_0 dark_weights_normed_gauss_ds_1_update_0_150(.clk(dark_weights_normed_gauss_ds_1_update_0_150_clk), .rst(dark_weights_normed_gauss_ds_1_update_0_150_rst), .start(dark_weights_normed_gauss_ds_1_update_0_150_start), .done(dark_weights_normed_gauss_ds_1_update_0_150_done), .src_in(dark_weights_normed_gauss_ds_1_update_0_150_src_in), .src_out(dark_weights_normed_gauss_ds_1_update_0_150_src_out), .out(dark_weights_normed_gauss_ds_1_update_0_150_out));
  assign dark_weights_normed_gauss_ds_1_update_0_150_clk = clk;
  assign dark_weights_normed_gauss_ds_1_update_0_150_rst = rst;
  assign dark_weights_normed_gauss_ds_1_update_0_150_start = start;
  // Bindings to dark_weights_normed_gauss_ds_1_update_0_150
    // dark_weights_normed_gauss_ds_1_update_0
  assign dark_weights_normed_gauss_ds_1_update_0 = dark_weights_normed_gauss_ds_1_update_0_150_out;

  // bright_weights_normed_gauss_blur_1_update_0_138
  logic [0:0] bright_weights_normed_gauss_blur_1_update_0_138_clk;
  logic [0:0] bright_weights_normed_gauss_blur_1_update_0_138_rst;
  logic [0:0] bright_weights_normed_gauss_blur_1_update_0_138_start;
  logic [0:0] bright_weights_normed_gauss_blur_1_update_0_138_done;
  logic [31:0] bright_weights_normed_gauss_blur_1_update_0_138_src_in;
  logic [31:0] bright_weights_normed_gauss_blur_1_update_0_138_src_out;
  logic [31:0] bright_weights_normed_gauss_blur_1_update_0_138_out;
  bright_weights_normed_gauss_blur_1_update_0 bright_weights_normed_gauss_blur_1_update_0_138(.clk(bright_weights_normed_gauss_blur_1_update_0_138_clk), .rst(bright_weights_normed_gauss_blur_1_update_0_138_rst), .start(bright_weights_normed_gauss_blur_1_update_0_138_start), .done(bright_weights_normed_gauss_blur_1_update_0_138_done), .src_in(bright_weights_normed_gauss_blur_1_update_0_138_src_in), .src_out(bright_weights_normed_gauss_blur_1_update_0_138_src_out), .out(bright_weights_normed_gauss_blur_1_update_0_138_out));
  assign bright_weights_normed_gauss_blur_1_update_0_138_clk = clk;
  assign bright_weights_normed_gauss_blur_1_update_0_138_rst = rst;
  assign bright_weights_normed_gauss_blur_1_update_0_138_start = start;
  // Bindings to bright_weights_normed_gauss_blur_1_update_0_138
    // bright_weights_normed_gauss_blur_1_update_0
  assign bright_weights_normed_gauss_blur_1_update_0 = bright_weights_normed_gauss_blur_1_update_0_138_out;

  // final_merged_2_update_0_141
  logic [0:0] final_merged_2_update_0_141_clk;
  logic [0:0] final_merged_2_update_0_141_rst;
  logic [0:0] final_merged_2_update_0_141_start;
  logic [0:0] final_merged_2_update_0_141_done;
  logic [31:0] final_merged_2_update_0_141_src_in;
  logic [31:0] final_merged_2_update_0_141_src_out;
  logic [31:0] final_merged_2_update_0_141_out;
  final_merged_2_update_0 final_merged_2_update_0_141(.clk(final_merged_2_update_0_141_clk), .rst(final_merged_2_update_0_141_rst), .start(final_merged_2_update_0_141_start), .done(final_merged_2_update_0_141_done), .src_in(final_merged_2_update_0_141_src_in), .src_out(final_merged_2_update_0_141_src_out), .out(final_merged_2_update_0_141_out));
  assign final_merged_2_update_0_141_clk = clk;
  assign final_merged_2_update_0_141_rst = rst;
  assign final_merged_2_update_0_141_start = start;
  // Bindings to final_merged_2_update_0_141
    // final_merged_2_update_0
  assign final_merged_2_update_0 = final_merged_2_update_0_141_out;

  // bright_weights_normed_gauss_blur_2_update_0_173
  logic [0:0] bright_weights_normed_gauss_blur_2_update_0_173_clk;
  logic [0:0] bright_weights_normed_gauss_blur_2_update_0_173_rst;
  logic [0:0] bright_weights_normed_gauss_blur_2_update_0_173_start;
  logic [0:0] bright_weights_normed_gauss_blur_2_update_0_173_done;
  logic [31:0] bright_weights_normed_gauss_blur_2_update_0_173_out;
  logic [31:0] bright_weights_normed_gauss_blur_2_update_0_173_src_in;
  logic [31:0] bright_weights_normed_gauss_blur_2_update_0_173_src_out;
  bright_weights_normed_gauss_blur_2_update_0 bright_weights_normed_gauss_blur_2_update_0_173(.clk(bright_weights_normed_gauss_blur_2_update_0_173_clk), .rst(bright_weights_normed_gauss_blur_2_update_0_173_rst), .start(bright_weights_normed_gauss_blur_2_update_0_173_start), .done(bright_weights_normed_gauss_blur_2_update_0_173_done), .out(bright_weights_normed_gauss_blur_2_update_0_173_out), .src_in(bright_weights_normed_gauss_blur_2_update_0_173_src_in), .src_out(bright_weights_normed_gauss_blur_2_update_0_173_src_out));
  assign bright_weights_normed_gauss_blur_2_update_0_173_clk = clk;
  assign bright_weights_normed_gauss_blur_2_update_0_173_rst = rst;
  assign bright_weights_normed_gauss_blur_2_update_0_173_start = start;
  // Bindings to bright_weights_normed_gauss_blur_2_update_0_173
    // bright_weights_normed_gauss_blur_2_update_0
  assign bright_weights_normed_gauss_blur_2_update_0 = bright_weights_normed_gauss_blur_2_update_0_173_out;

  // bright_laplace_diff_0_update_0_148
  logic [0:0] bright_laplace_diff_0_update_0_148_clk;
  logic [0:0] bright_laplace_diff_0_update_0_148_rst;
  logic [0:0] bright_laplace_diff_0_update_0_148_start;
  logic [0:0] bright_laplace_diff_0_update_0_148_done;
  logic [31:0] bright_laplace_diff_0_update_0_148_src_in;
  logic [31:0] bright_laplace_diff_0_update_0_148_src_out;
  logic [31:0] bright_laplace_diff_0_update_0_148_out;
  bright_laplace_diff_0_update_0 bright_laplace_diff_0_update_0_148(.clk(bright_laplace_diff_0_update_0_148_clk), .rst(bright_laplace_diff_0_update_0_148_rst), .start(bright_laplace_diff_0_update_0_148_start), .done(bright_laplace_diff_0_update_0_148_done), .src_in(bright_laplace_diff_0_update_0_148_src_in), .src_out(bright_laplace_diff_0_update_0_148_src_out), .out(bright_laplace_diff_0_update_0_148_out));
  assign bright_laplace_diff_0_update_0_148_clk = clk;
  assign bright_laplace_diff_0_update_0_148_rst = rst;
  assign bright_laplace_diff_0_update_0_148_start = start;
  // Bindings to bright_laplace_diff_0_update_0_148
    // bright_laplace_diff_0_update_0
  assign bright_laplace_diff_0_update_0 = bright_laplace_diff_0_update_0_148_out;

  // dark_gauss_ds_3_update_0_174
  logic [0:0] dark_gauss_ds_3_update_0_174_clk;
  logic [0:0] dark_gauss_ds_3_update_0_174_rst;
  logic [0:0] dark_gauss_ds_3_update_0_174_start;
  logic [0:0] dark_gauss_ds_3_update_0_174_done;
  logic [31:0] dark_gauss_ds_3_update_0_174_out;
  logic [31:0] dark_gauss_ds_3_update_0_174_src_in;
  logic [31:0] dark_gauss_ds_3_update_0_174_src_out;
  dark_gauss_ds_3_update_0 dark_gauss_ds_3_update_0_174(.clk(dark_gauss_ds_3_update_0_174_clk), .rst(dark_gauss_ds_3_update_0_174_rst), .start(dark_gauss_ds_3_update_0_174_start), .done(dark_gauss_ds_3_update_0_174_done), .out(dark_gauss_ds_3_update_0_174_out), .src_in(dark_gauss_ds_3_update_0_174_src_in), .src_out(dark_gauss_ds_3_update_0_174_src_out));
  assign dark_gauss_ds_3_update_0_174_clk = clk;
  assign dark_gauss_ds_3_update_0_174_rst = rst;
  assign dark_gauss_ds_3_update_0_174_start = start;
  // Bindings to dark_gauss_ds_3_update_0_174
    // dark_gauss_ds_3_update_0
  assign dark_gauss_ds_3_update_0 = dark_gauss_ds_3_update_0_174_out;

  // bright_weights_normed_gauss_ds_2_update_0_175
  logic [0:0] bright_weights_normed_gauss_ds_2_update_0_175_clk;
  logic [0:0] bright_weights_normed_gauss_ds_2_update_0_175_rst;
  logic [0:0] bright_weights_normed_gauss_ds_2_update_0_175_start;
  logic [0:0] bright_weights_normed_gauss_ds_2_update_0_175_done;
  logic [31:0] bright_weights_normed_gauss_ds_2_update_0_175_out;
  logic [31:0] bright_weights_normed_gauss_ds_2_update_0_175_src_in;
  logic [31:0] bright_weights_normed_gauss_ds_2_update_0_175_src_out;
  bright_weights_normed_gauss_ds_2_update_0 bright_weights_normed_gauss_ds_2_update_0_175(.clk(bright_weights_normed_gauss_ds_2_update_0_175_clk), .rst(bright_weights_normed_gauss_ds_2_update_0_175_rst), .start(bright_weights_normed_gauss_ds_2_update_0_175_start), .done(bright_weights_normed_gauss_ds_2_update_0_175_done), .out(bright_weights_normed_gauss_ds_2_update_0_175_out), .src_in(bright_weights_normed_gauss_ds_2_update_0_175_src_in), .src_out(bright_weights_normed_gauss_ds_2_update_0_175_src_out));
  assign bright_weights_normed_gauss_ds_2_update_0_175_clk = clk;
  assign bright_weights_normed_gauss_ds_2_update_0_175_rst = rst;
  assign bright_weights_normed_gauss_ds_2_update_0_175_start = start;
  // Bindings to bright_weights_normed_gauss_ds_2_update_0_175
    // bright_weights_normed_gauss_ds_2_update_0
  assign bright_weights_normed_gauss_ds_2_update_0 = bright_weights_normed_gauss_ds_2_update_0_175_out;

  // buf_bright_weights
  logic [0:0] buf_bright_weights_clk;
  logic [0:0] buf_bright_weights_rst;
  logic [0:0] buf_bright_weights_start;
  logic [0:0] buf_bright_weights_done;
  logic [0:0] buf_bright_weights_bright_weights_update_0_write_wen;
  logic [31:0] buf_bright_weights_weight_sums_update_0_read_dummy;
  logic [31:0] buf_bright_weights_bright_weights_update_0_write_wdata;
  logic [31:0] buf_bright_weights_bright_weights_normed_update_0_read_dummy;
  logic [31:0] buf_bright_weights_bright_weights_normed_update_0_read_rdata;
  logic [31:0] buf_bright_weights_weight_sums_update_0_read_rdata;
  bright_weights buf_bright_weights(.clk(buf_bright_weights_clk), .rst(buf_bright_weights_rst), .start(buf_bright_weights_start), .done(buf_bright_weights_done), .bright_weights_update_0_write_wen(buf_bright_weights_bright_weights_update_0_write_wen), .weight_sums_update_0_read_dummy(buf_bright_weights_weight_sums_update_0_read_dummy), .bright_weights_update_0_write_wdata(buf_bright_weights_bright_weights_update_0_write_wdata), .bright_weights_normed_update_0_read_dummy(buf_bright_weights_bright_weights_normed_update_0_read_dummy), .bright_weights_normed_update_0_read_rdata(buf_bright_weights_bright_weights_normed_update_0_read_rdata), .weight_sums_update_0_read_rdata(buf_bright_weights_weight_sums_update_0_read_rdata));
  assign buf_bright_weights_clk = clk;
  assign buf_bright_weights_rst = rst;
  assign buf_bright_weights_start = start;
  // Bindings to buf_bright_weights
    // bright_weights_bright_weights_update_0_write_write_5
  assign bright_weights_bright_weights_update_0_write_write_5 = buf_bright_weights_bright_weights_update_0_write_wdata;
  assign buf_bright_weights_bright_weights_update_0_write_wen = stage_8_active;
    // bright_weights_weight_sums_update_0_read_read_23
  assign bright_weights_weight_sums_update_0_read_read_23 = buf_bright_weights_weight_sums_update_0_read_rdata;
    // bright_weights_bright_weights_normed_update_0_read_read_48
  assign bright_weights_bright_weights_normed_update_0_read_read_48 = buf_bright_weights_bright_weights_normed_update_0_read_rdata;

  // buf_bright_laplace_diff_2
  logic [0:0] buf_bright_laplace_diff_2_clk;
  logic [0:0] buf_bright_laplace_diff_2_rst;
  logic [0:0] buf_bright_laplace_diff_2_start;
  logic [0:0] buf_bright_laplace_diff_2_done;
  logic [31:0] buf_bright_laplace_diff_2_fused_level_2_update_0_read_dummy;
  logic [0:0] buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wen;
  logic [31:0] buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_diff_2_fused_level_2_update_0_read_rdata;
  bright_laplace_diff_2 buf_bright_laplace_diff_2(.clk(buf_bright_laplace_diff_2_clk), .rst(buf_bright_laplace_diff_2_rst), .start(buf_bright_laplace_diff_2_start), .done(buf_bright_laplace_diff_2_done), .fused_level_2_update_0_read_dummy(buf_bright_laplace_diff_2_fused_level_2_update_0_read_dummy), .bright_laplace_diff_2_update_0_write_wen(buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wen), .bright_laplace_diff_2_update_0_write_wdata(buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wdata), .fused_level_2_update_0_read_rdata(buf_bright_laplace_diff_2_fused_level_2_update_0_read_rdata));
  assign buf_bright_laplace_diff_2_clk = clk;
  assign buf_bright_laplace_diff_2_rst = rst;
  assign buf_bright_laplace_diff_2_start = start;
  // Bindings to buf_bright_laplace_diff_2
    // bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84
  assign bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_write_84 = buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wdata;
  assign buf_bright_laplace_diff_2_bright_laplace_diff_2_update_0_write_wen = stage_121_active;
    // bright_laplace_diff_2_fused_level_2_update_0_read_read_107
  assign bright_laplace_diff_2_fused_level_2_update_0_read_read_107 = buf_bright_laplace_diff_2_fused_level_2_update_0_read_rdata;

  // buf_bright_laplace_us_0
  logic [0:0] buf_bright_laplace_us_0_clk;
  logic [0:0] buf_bright_laplace_us_0_rst;
  logic [0:0] buf_bright_laplace_us_0_start;
  logic [0:0] buf_bright_laplace_us_0_done;
  logic [0:0] buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wen;
  logic [31:0] buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_us_0_bright_laplace_diff_0_update_0_read_dummy;
  logic [31:0] buf_bright_laplace_us_0_bright_laplace_diff_0_update_0_read_rdata;
  bright_laplace_us_0 buf_bright_laplace_us_0(.clk(buf_bright_laplace_us_0_clk), .rst(buf_bright_laplace_us_0_rst), .start(buf_bright_laplace_us_0_start), .done(buf_bright_laplace_us_0_done), .bright_laplace_us_0_update_0_write_wen(buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wen), .bright_laplace_us_0_update_0_write_wdata(buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wdata), .bright_laplace_diff_0_update_0_read_dummy(buf_bright_laplace_us_0_bright_laplace_diff_0_update_0_read_dummy), .bright_laplace_diff_0_update_0_read_rdata(buf_bright_laplace_us_0_bright_laplace_diff_0_update_0_read_rdata));
  assign buf_bright_laplace_us_0_clk = clk;
  assign buf_bright_laplace_us_0_rst = rst;
  assign buf_bright_laplace_us_0_start = start;
  // Bindings to buf_bright_laplace_us_0
    // bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43
  assign bright_laplace_us_0_bright_laplace_diff_0_update_0_read_read_43 = buf_bright_laplace_us_0_bright_laplace_diff_0_update_0_read_rdata;
    // bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31
  assign bright_laplace_us_0_bright_laplace_us_0_update_0_write_write_31 = buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wdata;
  assign buf_bright_laplace_us_0_bright_laplace_us_0_update_0_write_wen = stage_46_active;

  // buf_bright_laplace_us_1
  logic [0:0] buf_bright_laplace_us_1_clk;
  logic [0:0] buf_bright_laplace_us_1_rst;
  logic [0:0] buf_bright_laplace_us_1_start;
  logic [0:0] buf_bright_laplace_us_1_done;
  logic [0:0] buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wen;
  logic [31:0] buf_bright_laplace_us_1_bright_laplace_diff_1_update_0_read_rdata;
  logic [31:0] buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_us_1_bright_laplace_diff_1_update_0_read_dummy;
  bright_laplace_us_1 buf_bright_laplace_us_1(.clk(buf_bright_laplace_us_1_clk), .rst(buf_bright_laplace_us_1_rst), .start(buf_bright_laplace_us_1_start), .done(buf_bright_laplace_us_1_done), .bright_laplace_us_1_update_0_write_wen(buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wen), .bright_laplace_diff_1_update_0_read_rdata(buf_bright_laplace_us_1_bright_laplace_diff_1_update_0_read_rdata), .bright_laplace_us_1_update_0_write_wdata(buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wdata), .bright_laplace_diff_1_update_0_read_dummy(buf_bright_laplace_us_1_bright_laplace_diff_1_update_0_read_dummy));
  assign buf_bright_laplace_us_1_clk = clk;
  assign buf_bright_laplace_us_1_rst = rst;
  assign buf_bright_laplace_us_1_start = start;
  // Bindings to buf_bright_laplace_us_1
    // bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41
  assign bright_laplace_us_1_bright_laplace_us_1_update_0_write_write_41 = buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wdata;
  assign buf_bright_laplace_us_1_bright_laplace_us_1_update_0_write_wen = stage_61_active;
    // bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68
  assign bright_laplace_us_1_bright_laplace_diff_1_update_0_read_read_68 = buf_bright_laplace_us_1_bright_laplace_diff_1_update_0_read_rdata;

  // buf_bright_laplace_us_2
  logic [0:0] buf_bright_laplace_us_2_clk;
  logic [0:0] buf_bright_laplace_us_2_rst;
  logic [0:0] buf_bright_laplace_us_2_start;
  logic [0:0] buf_bright_laplace_us_2_done;
  logic [0:0] buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wen;
  logic [31:0] buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wdata;
  logic [31:0] buf_bright_laplace_us_2_bright_laplace_diff_2_update_0_read_dummy;
  logic [31:0] buf_bright_laplace_us_2_bright_laplace_diff_2_update_0_read_rdata;
  bright_laplace_us_2 buf_bright_laplace_us_2(.clk(buf_bright_laplace_us_2_clk), .rst(buf_bright_laplace_us_2_rst), .start(buf_bright_laplace_us_2_start), .done(buf_bright_laplace_us_2_done), .bright_laplace_us_2_update_0_write_wen(buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wen), .bright_laplace_us_2_update_0_write_wdata(buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wdata), .bright_laplace_diff_2_update_0_read_dummy(buf_bright_laplace_us_2_bright_laplace_diff_2_update_0_read_dummy), .bright_laplace_diff_2_update_0_read_rdata(buf_bright_laplace_us_2_bright_laplace_diff_2_update_0_read_rdata));
  assign buf_bright_laplace_us_2_clk = clk;
  assign buf_bright_laplace_us_2_rst = rst;
  assign buf_bright_laplace_us_2_start = start;
  // Bindings to buf_bright_laplace_us_2
    // bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60
  assign bright_laplace_us_2_bright_laplace_us_2_update_0_write_write_60 = buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wdata;
  assign buf_bright_laplace_us_2_bright_laplace_us_2_update_0_write_wen = stage_88_active;
    // bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83
  assign bright_laplace_us_2_bright_laplace_diff_2_update_0_read_read_83 = buf_bright_laplace_us_2_bright_laplace_diff_2_update_0_read_rdata;

  // buf_dark
  logic [0:0] buf_dark_clk;
  logic [0:0] buf_dark_rst;
  logic [0:0] buf_dark_start;
  logic [0:0] buf_dark_done;
  logic [31:0] buf_dark_dark_update_0_write_wdata;
  logic [31:0] buf_dark_dark_weights_update_0_read_rdata;
  logic [31:0] buf_dark_dark_laplace_diff_0_update_0_read_rdata;
  logic [287:0] buf_dark_dark_gauss_blur_1_update_0_read_rdata;
  logic [31:0] buf_dark_dark_laplace_diff_0_update_0_read_dummy;
  logic [31:0] buf_dark_dark_weights_update_0_read_dummy;
  logic [287:0] buf_dark_dark_gauss_blur_1_update_0_read_dummy;
  logic [0:0] buf_dark_dark_update_0_write_wen;
  dark buf_dark(.clk(buf_dark_clk), .rst(buf_dark_rst), .start(buf_dark_start), .done(buf_dark_done), .dark_update_0_write_wdata(buf_dark_dark_update_0_write_wdata), .dark_weights_update_0_read_rdata(buf_dark_dark_weights_update_0_read_rdata), .dark_laplace_diff_0_update_0_read_rdata(buf_dark_dark_laplace_diff_0_update_0_read_rdata), .dark_gauss_blur_1_update_0_read_rdata(buf_dark_dark_gauss_blur_1_update_0_read_rdata), .dark_laplace_diff_0_update_0_read_dummy(buf_dark_dark_laplace_diff_0_update_0_read_dummy), .dark_weights_update_0_read_dummy(buf_dark_dark_weights_update_0_read_dummy), .dark_gauss_blur_1_update_0_read_dummy(buf_dark_dark_gauss_blur_1_update_0_read_dummy), .dark_update_0_write_wen(buf_dark_dark_update_0_write_wen));
  assign buf_dark_clk = clk;
  assign buf_dark_rst = rst;
  assign buf_dark_start = start;
  // Bindings to buf_dark
    // dark_dark_weights_update_0_read_read_8
  assign dark_dark_weights_update_0_read_read_8 = buf_dark_dark_weights_update_0_read_rdata;
    // dark_dark_update_0_write_write_7
  assign dark_dark_update_0_write_write_7 = buf_dark_dark_update_0_write_wdata;
  assign buf_dark_dark_update_0_write_wen = stage_11_active;
    // dark_dark_gauss_blur_1_update_0_read_read_10
  assign dark_dark_gauss_blur_1_update_0_read_read_10 = buf_dark_dark_gauss_blur_1_update_0_read_rdata;
    // dark_dark_laplace_diff_0_update_0_read_read_27
  assign dark_dark_laplace_diff_0_update_0_read_read_27 = buf_dark_dark_laplace_diff_0_update_0_read_rdata;

  // buf_bright_weights_normed
  logic [0:0] buf_bright_weights_normed_clk;
  logic [0:0] buf_bright_weights_normed_rst;
  logic [0:0] buf_bright_weights_normed_start;
  logic [0:0] buf_bright_weights_normed_done;
  logic [31:0] buf_bright_weights_normed_fused_level_0_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_fused_level_0_update_0_read_rdata;
  logic [0:0] buf_bright_weights_normed_bright_weights_normed_update_0_write_wen;
  logic [31:0] buf_bright_weights_normed_bright_weights_normed_update_0_write_wdata;
  logic [287:0] buf_bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_dummy;
  logic [287:0] buf_bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_rdata;
  bright_weights_normed buf_bright_weights_normed(.clk(buf_bright_weights_normed_clk), .rst(buf_bright_weights_normed_rst), .start(buf_bright_weights_normed_start), .done(buf_bright_weights_normed_done), .fused_level_0_update_0_read_dummy(buf_bright_weights_normed_fused_level_0_update_0_read_dummy), .fused_level_0_update_0_read_rdata(buf_bright_weights_normed_fused_level_0_update_0_read_rdata), .bright_weights_normed_update_0_write_wen(buf_bright_weights_normed_bright_weights_normed_update_0_write_wen), .bright_weights_normed_update_0_write_wdata(buf_bright_weights_normed_bright_weights_normed_update_0_write_wdata), .bright_weights_normed_gauss_blur_1_update_0_read_dummy(buf_bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_dummy), .bright_weights_normed_gauss_blur_1_update_0_read_rdata(buf_bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_rdata));
  assign buf_bright_weights_normed_clk = clk;
  assign buf_bright_weights_normed_rst = rst;
  assign buf_bright_weights_normed_start = start;
  // Bindings to buf_bright_weights_normed
    // bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55
  assign bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_read_55 = buf_bright_weights_normed_bright_weights_normed_gauss_blur_1_update_0_read_rdata;
    // bright_weights_normed_bright_weights_normed_update_0_write_write_50
  assign bright_weights_normed_bright_weights_normed_update_0_write_write_50 = buf_bright_weights_normed_bright_weights_normed_update_0_write_wdata;
  assign buf_bright_weights_normed_bright_weights_normed_update_0_write_wen = stage_73_active;
    // bright_weights_normed_fused_level_0_update_0_read_read_79
  assign bright_weights_normed_fused_level_0_update_0_read_read_79 = buf_bright_weights_normed_fused_level_0_update_0_read_rdata;

  // buf_dark_gauss_blur_1
  logic [0:0] buf_dark_gauss_blur_1_clk;
  logic [0:0] buf_dark_gauss_blur_1_rst;
  logic [0:0] buf_dark_gauss_blur_1_start;
  logic [0:0] buf_dark_gauss_blur_1_done;
  logic [0:0] buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wen;
  logic [31:0] buf_dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wdata;
  logic [31:0] buf_dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_rdata;
  dark_gauss_blur_1 buf_dark_gauss_blur_1(.clk(buf_dark_gauss_blur_1_clk), .rst(buf_dark_gauss_blur_1_rst), .start(buf_dark_gauss_blur_1_start), .done(buf_dark_gauss_blur_1_done), .dark_gauss_blur_1_update_0_write_wen(buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wen), .dark_gauss_ds_1_update_0_read_dummy(buf_dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_dummy), .dark_gauss_blur_1_update_0_write_wdata(buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wdata), .dark_gauss_ds_1_update_0_read_rdata(buf_dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_rdata));
  assign buf_dark_gauss_blur_1_clk = clk;
  assign buf_dark_gauss_blur_1_rst = rst;
  assign buf_dark_gauss_blur_1_start = start;
  // Bindings to buf_dark_gauss_blur_1
    // dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11
  assign dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_write_11 = buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wdata;
  assign buf_dark_gauss_blur_1_dark_gauss_blur_1_update_0_write_wen = stage_17_active;
    // dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14
  assign dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_read_14 = buf_dark_gauss_blur_1_dark_gauss_ds_1_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_blur_1
  logic [0:0] buf_bright_weights_normed_gauss_blur_1_clk;
  logic [0:0] buf_bright_weights_normed_gauss_blur_1_rst;
  logic [0:0] buf_bright_weights_normed_gauss_blur_1_start;
  logic [0:0] buf_bright_weights_normed_gauss_blur_1_done;
  logic [31:0] buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wdata;
  logic [0:0] buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wen;
  logic [31:0] buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_rdata;
  bright_weights_normed_gauss_blur_1 buf_bright_weights_normed_gauss_blur_1(.clk(buf_bright_weights_normed_gauss_blur_1_clk), .rst(buf_bright_weights_normed_gauss_blur_1_rst), .start(buf_bright_weights_normed_gauss_blur_1_start), .done(buf_bright_weights_normed_gauss_blur_1_done), .bright_weights_normed_gauss_blur_1_update_0_write_wdata(buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wdata), .bright_weights_normed_gauss_blur_1_update_0_write_wen(buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wen), .bright_weights_normed_gauss_ds_1_update_0_read_dummy(buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_dummy), .bright_weights_normed_gauss_ds_1_update_0_read_rdata(buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_rdata));
  assign buf_bright_weights_normed_gauss_blur_1_clk = clk;
  assign buf_bright_weights_normed_gauss_blur_1_rst = rst;
  assign buf_bright_weights_normed_gauss_blur_1_start = start;
  // Bindings to buf_bright_weights_normed_gauss_blur_1
    // bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_write_56 = buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_blur_1_update_0_write_wen = stage_82_active;
    // bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70
  assign bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_read_70 = buf_bright_weights_normed_gauss_blur_1_bright_weights_normed_gauss_ds_1_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_blur_2
  logic [0:0] buf_bright_weights_normed_gauss_blur_2_clk;
  logic [0:0] buf_bright_weights_normed_gauss_blur_2_rst;
  logic [0:0] buf_bright_weights_normed_gauss_blur_2_start;
  logic [0:0] buf_bright_weights_normed_gauss_blur_2_done;
  logic [0:0] buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wen;
  logic [31:0] buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wdata;
  logic [31:0] buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_rdata;
  bright_weights_normed_gauss_blur_2 buf_bright_weights_normed_gauss_blur_2(.clk(buf_bright_weights_normed_gauss_blur_2_clk), .rst(buf_bright_weights_normed_gauss_blur_2_rst), .start(buf_bright_weights_normed_gauss_blur_2_start), .done(buf_bright_weights_normed_gauss_blur_2_done), .bright_weights_normed_gauss_blur_2_update_0_write_wen(buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wen), .bright_weights_normed_gauss_blur_2_update_0_write_wdata(buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wdata), .bright_weights_normed_gauss_ds_2_update_0_read_dummy(buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_dummy), .bright_weights_normed_gauss_ds_2_update_0_read_rdata(buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_rdata));
  assign buf_bright_weights_normed_gauss_blur_2_clk = clk;
  assign buf_bright_weights_normed_gauss_blur_2_rst = rst;
  assign buf_bright_weights_normed_gauss_blur_2_start = start;
  // Bindings to buf_bright_weights_normed_gauss_blur_2
    // bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_write_91 = buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_blur_2_update_0_write_wen = stage_130_active;
    // bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96
  assign bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_read_96 = buf_bright_weights_normed_gauss_blur_2_bright_weights_normed_gauss_ds_2_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_blur_3
  logic [0:0] buf_bright_weights_normed_gauss_blur_3_clk;
  logic [0:0] buf_bright_weights_normed_gauss_blur_3_rst;
  logic [0:0] buf_bright_weights_normed_gauss_blur_3_start;
  logic [0:0] buf_bright_weights_normed_gauss_blur_3_done;
  logic [0:0] buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wen;
  logic [31:0] buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wdata;
  logic [31:0] buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_rdata;
  bright_weights_normed_gauss_blur_3 buf_bright_weights_normed_gauss_blur_3(.clk(buf_bright_weights_normed_gauss_blur_3_clk), .rst(buf_bright_weights_normed_gauss_blur_3_rst), .start(buf_bright_weights_normed_gauss_blur_3_start), .done(buf_bright_weights_normed_gauss_blur_3_done), .bright_weights_normed_gauss_blur_3_update_0_write_wen(buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wen), .bright_weights_normed_gauss_blur_3_update_0_write_wdata(buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wdata), .bright_weights_normed_gauss_ds_3_update_0_read_dummy(buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_dummy), .bright_weights_normed_gauss_ds_3_update_0_read_rdata(buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_rdata));
  assign buf_bright_weights_normed_gauss_blur_3_clk = clk;
  assign buf_bright_weights_normed_gauss_blur_3_rst = rst;
  assign buf_bright_weights_normed_gauss_blur_3_start = start;
  // Bindings to buf_bright_weights_normed_gauss_blur_3
    // bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_write_104 = buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_blur_3_update_0_write_wen = stage_149_active;
    // bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105
  assign bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_read_105 = buf_bright_weights_normed_gauss_blur_3_bright_weights_normed_gauss_ds_3_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_ds_1
  logic [0:0] buf_bright_weights_normed_gauss_ds_1_clk;
  logic [0:0] buf_bright_weights_normed_gauss_ds_1_rst;
  logic [0:0] buf_bright_weights_normed_gauss_ds_1_start;
  logic [0:0] buf_bright_weights_normed_gauss_ds_1_done;
  logic [287:0] buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_dummy;
  logic [0:0] buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wen;
  logic [31:0] buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wdata;
  logic [287:0] buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_rdata;
  logic [31:0] buf_bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata;
  bright_weights_normed_gauss_ds_1 buf_bright_weights_normed_gauss_ds_1(.clk(buf_bright_weights_normed_gauss_ds_1_clk), .rst(buf_bright_weights_normed_gauss_ds_1_rst), .start(buf_bright_weights_normed_gauss_ds_1_start), .done(buf_bright_weights_normed_gauss_ds_1_done), .bright_weights_normed_gauss_blur_2_update_0_read_dummy(buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_dummy), .bright_weights_normed_gauss_ds_1_update_0_write_wen(buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wen), .bright_weights_normed_gauss_ds_1_update_0_write_wdata(buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wdata), .bright_weights_normed_gauss_blur_2_update_0_read_rdata(buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_rdata), .fused_level_1_update_0_read_dummy(buf_bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_dummy), .fused_level_1_update_0_read_rdata(buf_bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata));
  assign buf_bright_weights_normed_gauss_ds_1_clk = clk;
  assign buf_bright_weights_normed_gauss_ds_1_rst = rst;
  assign buf_bright_weights_normed_gauss_ds_1_start = start;
  // Bindings to buf_bright_weights_normed_gauss_ds_1
    // bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_write_71 = buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_ds_1_update_0_write_wen = stage_104_active;
    // bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87
  assign bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_87 = buf_bright_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata;
    // bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90
  assign bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_read_90 = buf_bright_weights_normed_gauss_ds_1_bright_weights_normed_gauss_blur_2_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_ds_2
  logic [0:0] buf_bright_weights_normed_gauss_ds_2_clk;
  logic [0:0] buf_bright_weights_normed_gauss_ds_2_rst;
  logic [0:0] buf_bright_weights_normed_gauss_ds_2_start;
  logic [0:0] buf_bright_weights_normed_gauss_ds_2_done;
  logic [287:0] buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wdata;
  logic [0:0] buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wen;
  logic [287:0] buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_rdata;
  logic [31:0] buf_bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_dummy;
  logic [31:0] buf_bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata;
  bright_weights_normed_gauss_ds_2 buf_bright_weights_normed_gauss_ds_2(.clk(buf_bright_weights_normed_gauss_ds_2_clk), .rst(buf_bright_weights_normed_gauss_ds_2_rst), .start(buf_bright_weights_normed_gauss_ds_2_start), .done(buf_bright_weights_normed_gauss_ds_2_done), .bright_weights_normed_gauss_blur_3_update_0_read_dummy(buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_dummy), .bright_weights_normed_gauss_ds_2_update_0_write_wdata(buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wdata), .bright_weights_normed_gauss_ds_2_update_0_write_wen(buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wen), .bright_weights_normed_gauss_blur_3_update_0_read_rdata(buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_rdata), .fused_level_2_update_0_read_dummy(buf_bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_dummy), .fused_level_2_update_0_read_rdata(buf_bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata));
  assign buf_bright_weights_normed_gauss_ds_2_clk = clk;
  assign buf_bright_weights_normed_gauss_ds_2_rst = rst;
  assign buf_bright_weights_normed_gauss_ds_2_start = start;
  // Bindings to buf_bright_weights_normed_gauss_ds_2
    // bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_write_97 = buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_ds_2_update_0_write_wen = stage_139_active;
    // bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103
  assign bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_read_103 = buf_bright_weights_normed_gauss_ds_2_bright_weights_normed_gauss_blur_3_update_0_read_rdata;
    // bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109
  assign bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_109 = buf_bright_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata;

  // buf_bright_weights_normed_gauss_ds_3
  logic [0:0] buf_bright_weights_normed_gauss_ds_3_clk;
  logic [0:0] buf_bright_weights_normed_gauss_ds_3_rst;
  logic [0:0] buf_bright_weights_normed_gauss_ds_3_start;
  logic [0:0] buf_bright_weights_normed_gauss_ds_3_done;
  logic [31:0] buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wdata;
  logic [31:0] buf_bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata;
  logic [31:0] buf_bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_dummy;
  logic [0:0] buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wen;
  bright_weights_normed_gauss_ds_3 buf_bright_weights_normed_gauss_ds_3(.clk(buf_bright_weights_normed_gauss_ds_3_clk), .rst(buf_bright_weights_normed_gauss_ds_3_rst), .start(buf_bright_weights_normed_gauss_ds_3_start), .done(buf_bright_weights_normed_gauss_ds_3_done), .bright_weights_normed_gauss_ds_3_update_0_write_wdata(buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wdata), .fused_level_3_update_0_read_rdata(buf_bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata), .fused_level_3_update_0_read_dummy(buf_bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_dummy), .bright_weights_normed_gauss_ds_3_update_0_write_wen(buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wen));
  assign buf_bright_weights_normed_gauss_ds_3_clk = clk;
  assign buf_bright_weights_normed_gauss_ds_3_rst = rst;
  assign buf_bright_weights_normed_gauss_ds_3_start = start;
  // Bindings to buf_bright_weights_normed_gauss_ds_3
    // bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114
  assign bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_114 = buf_bright_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata;
    // bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106
  assign bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_write_106 = buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wdata;
  assign buf_bright_weights_normed_gauss_ds_3_bright_weights_normed_gauss_ds_3_update_0_write_wen = stage_152_active;

  // buf_dark_gauss_blur_2
  logic [0:0] buf_dark_gauss_blur_2_clk;
  logic [0:0] buf_dark_gauss_blur_2_rst;
  logic [0:0] buf_dark_gauss_blur_2_start;
  logic [0:0] buf_dark_gauss_blur_2_done;
  logic [31:0] buf_dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wdata;
  logic [0:0] buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wen;
  logic [31:0] buf_dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_dummy;
  dark_gauss_blur_2 buf_dark_gauss_blur_2(.clk(buf_dark_gauss_blur_2_clk), .rst(buf_dark_gauss_blur_2_rst), .start(buf_dark_gauss_blur_2_start), .done(buf_dark_gauss_blur_2_done), .dark_gauss_ds_2_update_0_read_rdata(buf_dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_rdata), .dark_gauss_blur_2_update_0_write_wdata(buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wdata), .dark_gauss_blur_2_update_0_write_wen(buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wen), .dark_gauss_ds_2_update_0_read_dummy(buf_dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_dummy));
  assign buf_dark_gauss_blur_2_clk = clk;
  assign buf_dark_gauss_blur_2_rst = rst;
  assign buf_dark_gauss_blur_2_start = start;
  // Bindings to buf_dark_gauss_blur_2
    // dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19
  assign dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_write_19 = buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wdata;
  assign buf_dark_gauss_blur_2_dark_gauss_blur_2_update_0_write_wen = stage_29_active;
    // dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34
  assign dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_read_34 = buf_dark_gauss_blur_2_dark_gauss_ds_2_update_0_read_rdata;

  // buf_dark_gauss_blur_3
  logic [0:0] buf_dark_gauss_blur_3_clk;
  logic [0:0] buf_dark_gauss_blur_3_rst;
  logic [0:0] buf_dark_gauss_blur_3_start;
  logic [0:0] buf_dark_gauss_blur_3_done;
  logic [0:0] buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wen;
  logic [31:0] buf_dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wdata;
  logic [31:0] buf_dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_rdata;
  dark_gauss_blur_3 buf_dark_gauss_blur_3(.clk(buf_dark_gauss_blur_3_clk), .rst(buf_dark_gauss_blur_3_rst), .start(buf_dark_gauss_blur_3_start), .done(buf_dark_gauss_blur_3_done), .dark_gauss_blur_3_update_0_write_wen(buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wen), .dark_gauss_ds_3_update_0_read_dummy(buf_dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_dummy), .dark_gauss_blur_3_update_0_write_wdata(buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wdata), .dark_gauss_ds_3_update_0_read_rdata(buf_dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_rdata));
  assign buf_dark_gauss_blur_3_clk = clk;
  assign buf_dark_gauss_blur_3_rst = rst;
  assign buf_dark_gauss_blur_3_start = start;
  // Bindings to buf_dark_gauss_blur_3
    // dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66
  assign dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_write_66 = buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wdata;
  assign buf_dark_gauss_blur_3_dark_gauss_blur_3_update_0_write_wen = stage_97_active;
    // dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92
  assign dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_read_92 = buf_dark_gauss_blur_3_dark_gauss_ds_3_update_0_read_rdata;

  // buf_dark_gauss_ds_1
  logic [0:0] buf_dark_gauss_ds_1_clk;
  logic [0:0] buf_dark_gauss_ds_1_rst;
  logic [0:0] buf_dark_gauss_ds_1_start;
  logic [0:0] buf_dark_gauss_ds_1_done;
  logic [287:0] buf_dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_1_dark_laplace_us_0_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_1_dark_laplace_us_0_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_dummy;
  logic [287:0] buf_dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_dummy;
  logic [0:0] buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wen;
  logic [31:0] buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wdata;
  dark_gauss_ds_1 buf_dark_gauss_ds_1(.clk(buf_dark_gauss_ds_1_clk), .rst(buf_dark_gauss_ds_1_rst), .start(buf_dark_gauss_ds_1_start), .done(buf_dark_gauss_ds_1_done), .dark_gauss_blur_2_update_0_read_rdata(buf_dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_rdata), .dark_laplace_us_0_update_0_read_rdata(buf_dark_gauss_ds_1_dark_laplace_us_0_update_0_read_rdata), .dark_laplace_us_0_update_0_read_dummy(buf_dark_gauss_ds_1_dark_laplace_us_0_update_0_read_dummy), .dark_laplace_diff_1_update_0_read_rdata(buf_dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_rdata), .dark_laplace_diff_1_update_0_read_dummy(buf_dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_dummy), .dark_gauss_blur_2_update_0_read_dummy(buf_dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_dummy), .dark_gauss_ds_1_update_0_write_wen(buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wen), .dark_gauss_ds_1_update_0_write_wdata(buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wdata));
  assign buf_dark_gauss_ds_1_clk = clk;
  assign buf_dark_gauss_ds_1_rst = rst;
  assign buf_dark_gauss_ds_1_start = start;
  // Bindings to buf_dark_gauss_ds_1
    // dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16
  assign dark_gauss_ds_1_dark_laplace_us_0_update_0_read_read_16 = buf_dark_gauss_ds_1_dark_laplace_us_0_update_0_read_rdata;
    // dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15
  assign dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_write_15 = buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wdata;
  assign buf_dark_gauss_ds_1_dark_gauss_ds_1_update_0_write_wen = stage_23_active;
    // dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18
  assign dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_read_18 = buf_dark_gauss_ds_1_dark_gauss_blur_2_update_0_read_rdata;
    // dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74
  assign dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_read_74 = buf_dark_gauss_ds_1_dark_laplace_diff_1_update_0_read_rdata;

  // buf_dark_gauss_ds_2
  logic [0:0] buf_dark_gauss_ds_2_clk;
  logic [0:0] buf_dark_gauss_ds_2_rst;
  logic [0:0] buf_dark_gauss_ds_2_start;
  logic [0:0] buf_dark_gauss_ds_2_done;
  logic [0:0] buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wen;
  logic [31:0] buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wdata;
  logic [287:0] buf_dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_dummy;
  logic [287:0] buf_dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_2_dark_laplace_us_1_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_ds_2_dark_laplace_us_1_update_0_read_rdata;
  dark_gauss_ds_2 buf_dark_gauss_ds_2(.clk(buf_dark_gauss_ds_2_clk), .rst(buf_dark_gauss_ds_2_rst), .start(buf_dark_gauss_ds_2_start), .done(buf_dark_gauss_ds_2_done), .dark_gauss_ds_2_update_0_write_wen(buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wen), .dark_gauss_ds_2_update_0_write_wdata(buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wdata), .dark_gauss_blur_3_update_0_read_dummy(buf_dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_dummy), .dark_gauss_blur_3_update_0_read_rdata(buf_dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_rdata), .dark_laplace_diff_2_update_0_read_dummy(buf_dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_dummy), .dark_laplace_diff_2_update_0_read_rdata(buf_dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_rdata), .dark_laplace_us_1_update_0_read_dummy(buf_dark_gauss_ds_2_dark_laplace_us_1_update_0_read_dummy), .dark_laplace_us_1_update_0_read_rdata(buf_dark_gauss_ds_2_dark_laplace_us_1_update_0_read_rdata));
  assign buf_dark_gauss_ds_2_clk = clk;
  assign buf_dark_gauss_ds_2_rst = rst;
  assign buf_dark_gauss_ds_2_start = start;
  // Bindings to buf_dark_gauss_ds_2
    // dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61
  assign dark_gauss_ds_2_dark_laplace_us_1_update_0_read_read_61 = buf_dark_gauss_ds_2_dark_laplace_us_1_update_0_read_rdata;
    // dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65
  assign dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_read_65 = buf_dark_gauss_ds_2_dark_gauss_blur_3_update_0_read_rdata;
    // dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35
  assign dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_write_35 = buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wdata;
  assign buf_dark_gauss_ds_2_dark_gauss_ds_2_update_0_write_wen = stage_52_active;
    // dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100
  assign dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_read_100 = buf_dark_gauss_ds_2_dark_laplace_diff_2_update_0_read_rdata;

  // buf_dark_gauss_ds_3
  logic [0:0] buf_dark_gauss_ds_3_clk;
  logic [0:0] buf_dark_gauss_ds_3_rst;
  logic [0:0] buf_dark_gauss_ds_3_start;
  logic [0:0] buf_dark_gauss_ds_3_done;
  logic [0:0] buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wen;
  logic [31:0] buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wdata;
  logic [31:0] buf_dark_gauss_ds_3_dark_laplace_us_2_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_ds_3_dark_laplace_us_2_update_0_read_rdata;
  logic [31:0] buf_dark_gauss_ds_3_fused_level_3_update_0_read_dummy;
  logic [31:0] buf_dark_gauss_ds_3_fused_level_3_update_0_read_rdata;
  dark_gauss_ds_3 buf_dark_gauss_ds_3(.clk(buf_dark_gauss_ds_3_clk), .rst(buf_dark_gauss_ds_3_rst), .start(buf_dark_gauss_ds_3_start), .done(buf_dark_gauss_ds_3_done), .dark_gauss_ds_3_update_0_write_wen(buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wen), .dark_gauss_ds_3_update_0_write_wdata(buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wdata), .dark_laplace_us_2_update_0_read_dummy(buf_dark_gauss_ds_3_dark_laplace_us_2_update_0_read_dummy), .dark_laplace_us_2_update_0_read_rdata(buf_dark_gauss_ds_3_dark_laplace_us_2_update_0_read_rdata), .fused_level_3_update_0_read_dummy(buf_dark_gauss_ds_3_fused_level_3_update_0_read_dummy), .fused_level_3_update_0_read_rdata(buf_dark_gauss_ds_3_fused_level_3_update_0_read_rdata));
  assign buf_dark_gauss_ds_3_clk = clk;
  assign buf_dark_gauss_ds_3_rst = rst;
  assign buf_dark_gauss_ds_3_start = start;
  // Bindings to buf_dark_gauss_ds_3
    // dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98
  assign dark_gauss_ds_3_dark_laplace_us_2_update_0_read_read_98 = buf_dark_gauss_ds_3_dark_laplace_us_2_update_0_read_rdata;
    // dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93
  assign dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_write_93 = buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wdata;
  assign buf_dark_gauss_ds_3_dark_gauss_ds_3_update_0_write_wen = stage_133_active;
    // dark_gauss_ds_3_fused_level_3_update_0_read_read_113
  assign dark_gauss_ds_3_fused_level_3_update_0_read_read_113 = buf_dark_gauss_ds_3_fused_level_3_update_0_read_rdata;

  // buf_dark_laplace_us_0
  logic [0:0] buf_dark_laplace_us_0_clk;
  logic [0:0] buf_dark_laplace_us_0_rst;
  logic [0:0] buf_dark_laplace_us_0_start;
  logic [0:0] buf_dark_laplace_us_0_done;
  logic [0:0] buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wen;
  logic [31:0] buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_us_0_dark_laplace_diff_0_update_0_read_dummy;
  logic [31:0] buf_dark_laplace_us_0_dark_laplace_diff_0_update_0_read_rdata;
  dark_laplace_us_0 buf_dark_laplace_us_0(.clk(buf_dark_laplace_us_0_clk), .rst(buf_dark_laplace_us_0_rst), .start(buf_dark_laplace_us_0_start), .done(buf_dark_laplace_us_0_done), .dark_laplace_us_0_update_0_write_wen(buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wen), .dark_laplace_us_0_update_0_write_wdata(buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wdata), .dark_laplace_diff_0_update_0_read_dummy(buf_dark_laplace_us_0_dark_laplace_diff_0_update_0_read_dummy), .dark_laplace_diff_0_update_0_read_rdata(buf_dark_laplace_us_0_dark_laplace_diff_0_update_0_read_rdata));
  assign buf_dark_laplace_us_0_clk = clk;
  assign buf_dark_laplace_us_0_rst = rst;
  assign buf_dark_laplace_us_0_start = start;
  // Bindings to buf_dark_laplace_us_0
    // dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17
  assign dark_laplace_us_0_dark_laplace_us_0_update_0_write_write_17 = buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wdata;
  assign buf_dark_laplace_us_0_dark_laplace_us_0_update_0_write_wen = stage_26_active;
    // dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28
  assign dark_laplace_us_0_dark_laplace_diff_0_update_0_read_read_28 = buf_dark_laplace_us_0_dark_laplace_diff_0_update_0_read_rdata;

  // buf_dark_laplace_diff_0
  logic [0:0] buf_dark_laplace_diff_0_clk;
  logic [0:0] buf_dark_laplace_diff_0_rst;
  logic [0:0] buf_dark_laplace_diff_0_start;
  logic [0:0] buf_dark_laplace_diff_0_done;
  logic [31:0] buf_dark_laplace_diff_0_fused_level_0_update_0_read_dummy;
  logic [0:0] buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wen;
  logic [31:0] buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_diff_0_fused_level_0_update_0_read_rdata;
  dark_laplace_diff_0 buf_dark_laplace_diff_0(.clk(buf_dark_laplace_diff_0_clk), .rst(buf_dark_laplace_diff_0_rst), .start(buf_dark_laplace_diff_0_start), .done(buf_dark_laplace_diff_0_done), .fused_level_0_update_0_read_dummy(buf_dark_laplace_diff_0_fused_level_0_update_0_read_dummy), .dark_laplace_diff_0_update_0_write_wen(buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wen), .dark_laplace_diff_0_update_0_write_wdata(buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wdata), .fused_level_0_update_0_read_rdata(buf_dark_laplace_diff_0_fused_level_0_update_0_read_rdata));
  assign buf_dark_laplace_diff_0_clk = clk;
  assign buf_dark_laplace_diff_0_rst = rst;
  assign buf_dark_laplace_diff_0_start = start;
  // Bindings to buf_dark_laplace_diff_0
    // dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29
  assign dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_write_29 = buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wdata;
  assign buf_dark_laplace_diff_0_dark_laplace_diff_0_update_0_write_wen = stage_43_active;
    // dark_laplace_diff_0_fused_level_0_update_0_read_read_78
  assign dark_laplace_diff_0_fused_level_0_update_0_read_read_78 = buf_dark_laplace_diff_0_fused_level_0_update_0_read_rdata;

  // buf_dark_laplace_diff_1
  logic [0:0] buf_dark_laplace_diff_1_clk;
  logic [0:0] buf_dark_laplace_diff_1_rst;
  logic [0:0] buf_dark_laplace_diff_1_start;
  logic [0:0] buf_dark_laplace_diff_1_done;
  logic [0:0] buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wen;
  logic [31:0] buf_dark_laplace_diff_1_fused_level_1_update_0_read_dummy;
  logic [31:0] buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_diff_1_fused_level_1_update_0_read_rdata;
  dark_laplace_diff_1 buf_dark_laplace_diff_1(.clk(buf_dark_laplace_diff_1_clk), .rst(buf_dark_laplace_diff_1_rst), .start(buf_dark_laplace_diff_1_start), .done(buf_dark_laplace_diff_1_done), .dark_laplace_diff_1_update_0_write_wen(buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wen), .fused_level_1_update_0_read_dummy(buf_dark_laplace_diff_1_fused_level_1_update_0_read_dummy), .dark_laplace_diff_1_update_0_write_wdata(buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wdata), .fused_level_1_update_0_read_rdata(buf_dark_laplace_diff_1_fused_level_1_update_0_read_rdata));
  assign buf_dark_laplace_diff_1_clk = clk;
  assign buf_dark_laplace_diff_1_rst = rst;
  assign buf_dark_laplace_diff_1_start = start;
  // Bindings to buf_dark_laplace_diff_1
    // dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76
  assign dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_write_76 = buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wdata;
  assign buf_dark_laplace_diff_1_dark_laplace_diff_1_update_0_write_wen = stage_111_active;
    // dark_laplace_diff_1_fused_level_1_update_0_read_read_86
  assign dark_laplace_diff_1_fused_level_1_update_0_read_read_86 = buf_dark_laplace_diff_1_fused_level_1_update_0_read_rdata;

  // buf_dark_laplace_diff_2
  logic [0:0] buf_dark_laplace_diff_2_clk;
  logic [0:0] buf_dark_laplace_diff_2_rst;
  logic [0:0] buf_dark_laplace_diff_2_start;
  logic [0:0] buf_dark_laplace_diff_2_done;
  logic [31:0] buf_dark_laplace_diff_2_fused_level_2_update_0_read_dummy;
  logic [0:0] buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wen;
  logic [31:0] buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_diff_2_fused_level_2_update_0_read_rdata;
  dark_laplace_diff_2 buf_dark_laplace_diff_2(.clk(buf_dark_laplace_diff_2_clk), .rst(buf_dark_laplace_diff_2_rst), .start(buf_dark_laplace_diff_2_start), .done(buf_dark_laplace_diff_2_done), .fused_level_2_update_0_read_dummy(buf_dark_laplace_diff_2_fused_level_2_update_0_read_dummy), .dark_laplace_diff_2_update_0_write_wen(buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wen), .dark_laplace_diff_2_update_0_write_wdata(buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wdata), .fused_level_2_update_0_read_rdata(buf_dark_laplace_diff_2_fused_level_2_update_0_read_rdata));
  assign buf_dark_laplace_diff_2_clk = clk;
  assign buf_dark_laplace_diff_2_rst = rst;
  assign buf_dark_laplace_diff_2_start = start;
  // Bindings to buf_dark_laplace_diff_2
    // dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102
  assign dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_write_102 = buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wdata;
  assign buf_dark_laplace_diff_2_dark_laplace_diff_2_update_0_write_wen = stage_146_active;
    // dark_laplace_diff_2_fused_level_2_update_0_read_read_108
  assign dark_laplace_diff_2_fused_level_2_update_0_read_read_108 = buf_dark_laplace_diff_2_fused_level_2_update_0_read_rdata;

  // buf_dark_laplace_us_1
  logic [0:0] buf_dark_laplace_us_1_clk;
  logic [0:0] buf_dark_laplace_us_1_rst;
  logic [0:0] buf_dark_laplace_us_1_start;
  logic [0:0] buf_dark_laplace_us_1_done;
  logic [0:0] buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wen;
  logic [31:0] buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_us_1_dark_laplace_diff_1_update_0_read_dummy;
  logic [31:0] buf_dark_laplace_us_1_dark_laplace_diff_1_update_0_read_rdata;
  dark_laplace_us_1 buf_dark_laplace_us_1(.clk(buf_dark_laplace_us_1_clk), .rst(buf_dark_laplace_us_1_rst), .start(buf_dark_laplace_us_1_start), .done(buf_dark_laplace_us_1_done), .dark_laplace_us_1_update_0_write_wen(buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wen), .dark_laplace_us_1_update_0_write_wdata(buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wdata), .dark_laplace_diff_1_update_0_read_dummy(buf_dark_laplace_us_1_dark_laplace_diff_1_update_0_read_dummy), .dark_laplace_diff_1_update_0_read_rdata(buf_dark_laplace_us_1_dark_laplace_diff_1_update_0_read_rdata));
  assign buf_dark_laplace_us_1_clk = clk;
  assign buf_dark_laplace_us_1_rst = rst;
  assign buf_dark_laplace_us_1_start = start;
  // Bindings to buf_dark_laplace_us_1
    // dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62
  assign dark_laplace_us_1_dark_laplace_us_1_update_0_write_write_62 = buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wdata;
  assign buf_dark_laplace_us_1_dark_laplace_us_1_update_0_write_wen = stage_91_active;
    // dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75
  assign dark_laplace_us_1_dark_laplace_diff_1_update_0_read_read_75 = buf_dark_laplace_us_1_dark_laplace_diff_1_update_0_read_rdata;

  // buf_dark_laplace_us_2
  logic [0:0] buf_dark_laplace_us_2_clk;
  logic [0:0] buf_dark_laplace_us_2_rst;
  logic [0:0] buf_dark_laplace_us_2_start;
  logic [0:0] buf_dark_laplace_us_2_done;
  logic [0:0] buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wen;
  logic [31:0] buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wdata;
  logic [31:0] buf_dark_laplace_us_2_dark_laplace_diff_2_update_0_read_dummy;
  logic [31:0] buf_dark_laplace_us_2_dark_laplace_diff_2_update_0_read_rdata;
  dark_laplace_us_2 buf_dark_laplace_us_2(.clk(buf_dark_laplace_us_2_clk), .rst(buf_dark_laplace_us_2_rst), .start(buf_dark_laplace_us_2_start), .done(buf_dark_laplace_us_2_done), .dark_laplace_us_2_update_0_write_wen(buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wen), .dark_laplace_us_2_update_0_write_wdata(buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wdata), .dark_laplace_diff_2_update_0_read_dummy(buf_dark_laplace_us_2_dark_laplace_diff_2_update_0_read_dummy), .dark_laplace_diff_2_update_0_read_rdata(buf_dark_laplace_us_2_dark_laplace_diff_2_update_0_read_rdata));
  assign buf_dark_laplace_us_2_clk = clk;
  assign buf_dark_laplace_us_2_rst = rst;
  assign buf_dark_laplace_us_2_start = start;
  // Bindings to buf_dark_laplace_us_2
    // dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99
  assign dark_laplace_us_2_dark_laplace_us_2_update_0_write_write_99 = buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wdata;
  assign buf_dark_laplace_us_2_dark_laplace_us_2_update_0_write_wen = stage_142_active;
    // dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101
  assign dark_laplace_us_2_dark_laplace_diff_2_update_0_read_read_101 = buf_dark_laplace_us_2_dark_laplace_diff_2_update_0_read_rdata;

  // buf_dark_weights
  logic [0:0] buf_dark_weights_clk;
  logic [0:0] buf_dark_weights_rst;
  logic [0:0] buf_dark_weights_start;
  logic [0:0] buf_dark_weights_done;
  logic [0:0] buf_dark_weights_dark_weights_update_0_write_wen;
  logic [31:0] buf_dark_weights_dark_weights_update_0_write_wdata;
  logic [31:0] buf_dark_weights_weight_sums_update_0_read_dummy;
  logic [31:0] buf_dark_weights_dark_weights_normed_update_0_read_dummy;
  logic [31:0] buf_dark_weights_dark_weights_normed_update_0_read_rdata;
  logic [31:0] buf_dark_weights_weight_sums_update_0_read_rdata;
  dark_weights buf_dark_weights(.clk(buf_dark_weights_clk), .rst(buf_dark_weights_rst), .start(buf_dark_weights_start), .done(buf_dark_weights_done), .dark_weights_update_0_write_wen(buf_dark_weights_dark_weights_update_0_write_wen), .dark_weights_update_0_write_wdata(buf_dark_weights_dark_weights_update_0_write_wdata), .weight_sums_update_0_read_dummy(buf_dark_weights_weight_sums_update_0_read_dummy), .dark_weights_normed_update_0_read_dummy(buf_dark_weights_dark_weights_normed_update_0_read_dummy), .dark_weights_normed_update_0_read_rdata(buf_dark_weights_dark_weights_normed_update_0_read_rdata), .weight_sums_update_0_read_rdata(buf_dark_weights_weight_sums_update_0_read_rdata));
  assign buf_dark_weights_clk = clk;
  assign buf_dark_weights_rst = rst;
  assign buf_dark_weights_start = start;
  // Bindings to buf_dark_weights
    // dark_weights_dark_weights_update_0_write_write_9
  assign dark_weights_dark_weights_update_0_write_write_9 = buf_dark_weights_dark_weights_update_0_write_wdata;
  assign buf_dark_weights_dark_weights_update_0_write_wen = stage_14_active;
    // dark_weights_weight_sums_update_0_read_read_22
  assign dark_weights_weight_sums_update_0_read_read_22 = buf_dark_weights_weight_sums_update_0_read_rdata;
    // dark_weights_dark_weights_normed_update_0_read_read_45
  assign dark_weights_dark_weights_normed_update_0_read_read_45 = buf_dark_weights_dark_weights_normed_update_0_read_rdata;

  // buf_dark_weights_normed_gauss_ds_1
  logic [0:0] buf_dark_weights_normed_gauss_ds_1_clk;
  logic [0:0] buf_dark_weights_normed_gauss_ds_1_rst;
  logic [0:0] buf_dark_weights_normed_gauss_ds_1_start;
  logic [0:0] buf_dark_weights_normed_gauss_ds_1_done;
  logic [31:0] buf_dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata;
  logic [31:0] buf_dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_dummy;
  logic [287:0] buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_rdata;
  logic [31:0] buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wdata;
  logic [0:0] buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wen;
  logic [287:0] buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_dummy;
  dark_weights_normed_gauss_ds_1 buf_dark_weights_normed_gauss_ds_1(.clk(buf_dark_weights_normed_gauss_ds_1_clk), .rst(buf_dark_weights_normed_gauss_ds_1_rst), .start(buf_dark_weights_normed_gauss_ds_1_start), .done(buf_dark_weights_normed_gauss_ds_1_done), .fused_level_1_update_0_read_rdata(buf_dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata), .fused_level_1_update_0_read_dummy(buf_dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_dummy), .dark_weights_normed_gauss_blur_2_update_0_read_rdata(buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_rdata), .dark_weights_normed_gauss_ds_1_update_0_write_wdata(buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wdata), .dark_weights_normed_gauss_ds_1_update_0_write_wen(buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wen), .dark_weights_normed_gauss_blur_2_update_0_read_dummy(buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_dummy));
  assign buf_dark_weights_normed_gauss_ds_1_clk = clk;
  assign buf_dark_weights_normed_gauss_ds_1_rst = rst;
  assign buf_dark_weights_normed_gauss_ds_1_start = start;
  // Bindings to buf_dark_weights_normed_gauss_ds_1
    // dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_read_57 = buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_blur_2_update_0_read_rdata;
    // dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54
  assign dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_write_54 = buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_ds_1_dark_weights_normed_gauss_ds_1_update_0_write_wen = stage_79_active;
    // dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88
  assign dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_read_88 = buf_dark_weights_normed_gauss_ds_1_fused_level_1_update_0_read_rdata;

  // buf_dark_weights_normed
  logic [0:0] buf_dark_weights_normed_clk;
  logic [0:0] buf_dark_weights_normed_rst;
  logic [0:0] buf_dark_weights_normed_start;
  logic [0:0] buf_dark_weights_normed_done;
  logic [31:0] buf_dark_weights_normed_fused_level_0_update_0_read_dummy;
  logic [0:0] buf_dark_weights_normed_dark_weights_normed_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_dark_weights_normed_update_0_write_wdata;
  logic [287:0] buf_dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_dummy;
  logic [287:0] buf_dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_rdata;
  logic [31:0] buf_dark_weights_normed_fused_level_0_update_0_read_rdata;
  dark_weights_normed buf_dark_weights_normed(.clk(buf_dark_weights_normed_clk), .rst(buf_dark_weights_normed_rst), .start(buf_dark_weights_normed_start), .done(buf_dark_weights_normed_done), .fused_level_0_update_0_read_dummy(buf_dark_weights_normed_fused_level_0_update_0_read_dummy), .dark_weights_normed_update_0_write_wen(buf_dark_weights_normed_dark_weights_normed_update_0_write_wen), .dark_weights_normed_update_0_write_wdata(buf_dark_weights_normed_dark_weights_normed_update_0_write_wdata), .dark_weights_normed_gauss_blur_1_update_0_read_dummy(buf_dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_dummy), .dark_weights_normed_gauss_blur_1_update_0_read_rdata(buf_dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_rdata), .fused_level_0_update_0_read_rdata(buf_dark_weights_normed_fused_level_0_update_0_read_rdata));
  assign buf_dark_weights_normed_clk = clk;
  assign buf_dark_weights_normed_rst = rst;
  assign buf_dark_weights_normed_start = start;
  // Bindings to buf_dark_weights_normed
    // dark_weights_normed_dark_weights_normed_update_0_write_write_47
  assign dark_weights_normed_dark_weights_normed_update_0_write_write_47 = buf_dark_weights_normed_dark_weights_normed_update_0_write_wdata;
  assign buf_dark_weights_normed_dark_weights_normed_update_0_write_wen = stage_69_active;
    // dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51
  assign dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_read_51 = buf_dark_weights_normed_dark_weights_normed_gauss_blur_1_update_0_read_rdata;
    // dark_weights_normed_fused_level_0_update_0_read_read_80
  assign dark_weights_normed_fused_level_0_update_0_read_read_80 = buf_dark_weights_normed_fused_level_0_update_0_read_rdata;

  // buf_dark_weights_normed_gauss_blur_1
  logic [0:0] buf_dark_weights_normed_gauss_blur_1_clk;
  logic [0:0] buf_dark_weights_normed_gauss_blur_1_rst;
  logic [0:0] buf_dark_weights_normed_gauss_blur_1_start;
  logic [0:0] buf_dark_weights_normed_gauss_blur_1_done;
  logic [31:0] buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wdata;
  logic [31:0] buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_dummy;
  logic [0:0] buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_rdata;
  dark_weights_normed_gauss_blur_1 buf_dark_weights_normed_gauss_blur_1(.clk(buf_dark_weights_normed_gauss_blur_1_clk), .rst(buf_dark_weights_normed_gauss_blur_1_rst), .start(buf_dark_weights_normed_gauss_blur_1_start), .done(buf_dark_weights_normed_gauss_blur_1_done), .dark_weights_normed_gauss_blur_1_update_0_write_wdata(buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wdata), .dark_weights_normed_gauss_ds_1_update_0_read_dummy(buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_dummy), .dark_weights_normed_gauss_blur_1_update_0_write_wen(buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wen), .dark_weights_normed_gauss_ds_1_update_0_read_rdata(buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_rdata));
  assign buf_dark_weights_normed_gauss_blur_1_clk = clk;
  assign buf_dark_weights_normed_gauss_blur_1_rst = rst;
  assign buf_dark_weights_normed_gauss_blur_1_start = start;
  // Bindings to buf_dark_weights_normed_gauss_blur_1
    // dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_read_53 = buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_ds_1_update_0_read_rdata;
    // dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52
  assign dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_write_52 = buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_blur_1_dark_weights_normed_gauss_blur_1_update_0_write_wen = stage_76_active;

  // buf_dark_weights_normed_gauss_blur_2
  logic [0:0] buf_dark_weights_normed_gauss_blur_2_clk;
  logic [0:0] buf_dark_weights_normed_gauss_blur_2_rst;
  logic [0:0] buf_dark_weights_normed_gauss_blur_2_start;
  logic [0:0] buf_dark_weights_normed_gauss_blur_2_done;
  logic [0:0] buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wdata;
  logic [31:0] buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_dummy;
  logic [31:0] buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_rdata;
  dark_weights_normed_gauss_blur_2 buf_dark_weights_normed_gauss_blur_2(.clk(buf_dark_weights_normed_gauss_blur_2_clk), .rst(buf_dark_weights_normed_gauss_blur_2_rst), .start(buf_dark_weights_normed_gauss_blur_2_start), .done(buf_dark_weights_normed_gauss_blur_2_done), .dark_weights_normed_gauss_blur_2_update_0_write_wen(buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wen), .dark_weights_normed_gauss_blur_2_update_0_write_wdata(buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wdata), .dark_weights_normed_gauss_ds_2_update_0_read_dummy(buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_dummy), .dark_weights_normed_gauss_ds_2_update_0_read_rdata(buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_rdata));
  assign buf_dark_weights_normed_gauss_blur_2_clk = clk;
  assign buf_dark_weights_normed_gauss_blur_2_rst = rst;
  assign buf_dark_weights_normed_gauss_blur_2_start = start;
  // Bindings to buf_dark_weights_normed_gauss_blur_2
    // dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_write_58 = buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_blur_2_update_0_write_wen = stage_85_active;
    // dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63
  assign dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_read_63 = buf_dark_weights_normed_gauss_blur_2_dark_weights_normed_gauss_ds_2_update_0_read_rdata;

  // buf_dark_weights_normed_gauss_blur_3
  logic [0:0] buf_dark_weights_normed_gauss_blur_3_clk;
  logic [0:0] buf_dark_weights_normed_gauss_blur_3_rst;
  logic [0:0] buf_dark_weights_normed_gauss_blur_3_start;
  logic [0:0] buf_dark_weights_normed_gauss_blur_3_done;
  logic [0:0] buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wdata;
  logic [31:0] buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_dummy;
  logic [31:0] buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_rdata;
  dark_weights_normed_gauss_blur_3 buf_dark_weights_normed_gauss_blur_3(.clk(buf_dark_weights_normed_gauss_blur_3_clk), .rst(buf_dark_weights_normed_gauss_blur_3_rst), .start(buf_dark_weights_normed_gauss_blur_3_start), .done(buf_dark_weights_normed_gauss_blur_3_done), .dark_weights_normed_gauss_blur_3_update_0_write_wen(buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wen), .dark_weights_normed_gauss_blur_3_update_0_write_wdata(buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wdata), .dark_weights_normed_gauss_ds_3_update_0_read_dummy(buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_dummy), .dark_weights_normed_gauss_ds_3_update_0_read_rdata(buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_rdata));
  assign buf_dark_weights_normed_gauss_blur_3_clk = clk;
  assign buf_dark_weights_normed_gauss_blur_3_rst = rst;
  assign buf_dark_weights_normed_gauss_blur_3_start = start;
  // Bindings to buf_dark_weights_normed_gauss_blur_3
    // dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_read_94 = buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_ds_3_update_0_read_rdata;
    // dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73
  assign dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_write_73 = buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_blur_3_dark_weights_normed_gauss_blur_3_update_0_write_wen = stage_107_active;

  // buf_final_merged_0
  logic [0:0] buf_final_merged_0_clk;
  logic [0:0] buf_final_merged_0_rst;
  logic [0:0] buf_final_merged_0_start;
  logic [0:0] buf_final_merged_0_done;
  logic [0:0] buf_final_merged_0_final_merged_0_update_0_write_wen;
  logic [31:0] buf_final_merged_0_final_merged_0_update_0_write_wdata;
  logic [31:0] buf_final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_dummy;
  logic [31:0] buf_final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_rdata;
  final_merged_0 buf_final_merged_0(.clk(buf_final_merged_0_clk), .rst(buf_final_merged_0_rst), .start(buf_final_merged_0_start), .done(buf_final_merged_0_done), .final_merged_0_update_0_write_wen(buf_final_merged_0_final_merged_0_update_0_write_wen), .final_merged_0_update_0_write_wdata(buf_final_merged_0_final_merged_0_update_0_write_wdata), .pyramid_synthetic_exposure_fusion_update_0_read_dummy(buf_final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_dummy), .pyramid_synthetic_exposure_fusion_update_0_read_rdata(buf_final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_rdata));
  assign buf_final_merged_0_clk = clk;
  assign buf_final_merged_0_rst = rst;
  assign buf_final_merged_0_start = start;
  // Bindings to buf_final_merged_0
    // final_merged_0_final_merged_0_update_0_write_write_125
  assign final_merged_0_final_merged_0_update_0_write_write_125 = buf_final_merged_0_final_merged_0_update_0_write_wdata;
  assign buf_final_merged_0_final_merged_0_update_0_write_wen = stage_176_active;
    // final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126
  assign final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_read_126 = buf_final_merged_0_pyramid_synthetic_exposure_fusion_update_0_read_rdata;

  // buf_dark_weights_normed_gauss_ds_2
  logic [0:0] buf_dark_weights_normed_gauss_ds_2_clk;
  logic [0:0] buf_dark_weights_normed_gauss_ds_2_rst;
  logic [0:0] buf_dark_weights_normed_gauss_ds_2_start;
  logic [0:0] buf_dark_weights_normed_gauss_ds_2_done;
  logic [31:0] buf_dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_dummy;
  logic [287:0] buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_dummy;
  logic [0:0] buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wdata;
  logic [287:0] buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_rdata;
  logic [31:0] buf_dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata;
  dark_weights_normed_gauss_ds_2 buf_dark_weights_normed_gauss_ds_2(.clk(buf_dark_weights_normed_gauss_ds_2_clk), .rst(buf_dark_weights_normed_gauss_ds_2_rst), .start(buf_dark_weights_normed_gauss_ds_2_start), .done(buf_dark_weights_normed_gauss_ds_2_done), .fused_level_2_update_0_read_dummy(buf_dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_dummy), .dark_weights_normed_gauss_blur_3_update_0_read_dummy(buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_dummy), .dark_weights_normed_gauss_ds_2_update_0_write_wen(buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wen), .dark_weights_normed_gauss_ds_2_update_0_write_wdata(buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wdata), .dark_weights_normed_gauss_blur_3_update_0_read_rdata(buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_rdata), .fused_level_2_update_0_read_rdata(buf_dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata));
  assign buf_dark_weights_normed_gauss_ds_2_clk = clk;
  assign buf_dark_weights_normed_gauss_ds_2_rst = rst;
  assign buf_dark_weights_normed_gauss_ds_2_start = start;
  // Bindings to buf_dark_weights_normed_gauss_ds_2
    // dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_read_72 = buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_blur_3_update_0_read_rdata;
    // dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64
  assign dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_write_64 = buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_ds_2_dark_weights_normed_gauss_ds_2_update_0_write_wen = stage_94_active;
    // dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110
  assign dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_read_110 = buf_dark_weights_normed_gauss_ds_2_fused_level_2_update_0_read_rdata;

  // buf_dark_weights_normed_gauss_ds_3
  logic [0:0] buf_dark_weights_normed_gauss_ds_3_clk;
  logic [0:0] buf_dark_weights_normed_gauss_ds_3_rst;
  logic [0:0] buf_dark_weights_normed_gauss_ds_3_start;
  logic [0:0] buf_dark_weights_normed_gauss_ds_3_done;
  logic [31:0] buf_dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_dummy;
  logic [0:0] buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wen;
  logic [31:0] buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wdata;
  logic [31:0] buf_dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata;
  dark_weights_normed_gauss_ds_3 buf_dark_weights_normed_gauss_ds_3(.clk(buf_dark_weights_normed_gauss_ds_3_clk), .rst(buf_dark_weights_normed_gauss_ds_3_rst), .start(buf_dark_weights_normed_gauss_ds_3_start), .done(buf_dark_weights_normed_gauss_ds_3_done), .fused_level_3_update_0_read_dummy(buf_dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_dummy), .dark_weights_normed_gauss_ds_3_update_0_write_wen(buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wen), .dark_weights_normed_gauss_ds_3_update_0_write_wdata(buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wdata), .fused_level_3_update_0_read_rdata(buf_dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata));
  assign buf_dark_weights_normed_gauss_ds_3_clk = clk;
  assign buf_dark_weights_normed_gauss_ds_3_rst = rst;
  assign buf_dark_weights_normed_gauss_ds_3_start = start;
  // Bindings to buf_dark_weights_normed_gauss_ds_3
    // dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115
  assign dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_read_115 = buf_dark_weights_normed_gauss_ds_3_fused_level_3_update_0_read_rdata;
    // dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95
  assign dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_write_95 = buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wdata;
  assign buf_dark_weights_normed_gauss_ds_3_dark_weights_normed_gauss_ds_3_update_0_write_wen = stage_136_active;

  // buf_final_merged_1
  logic [0:0] buf_final_merged_1_clk;
  logic [0:0] buf_final_merged_1_rst;
  logic [0:0] buf_final_merged_1_start;
  logic [0:0] buf_final_merged_1_done;
  logic [0:0] buf_final_merged_1_final_merged_1_update_0_write_wen;
  logic [31:0] buf_final_merged_1_final_merged_1_update_0_write_wdata;
  logic [31:0] buf_final_merged_1_final_merged_0_update_0_read_dummy;
  logic [31:0] buf_final_merged_1_final_merged_0_update_0_read_rdata;
  final_merged_1 buf_final_merged_1(.clk(buf_final_merged_1_clk), .rst(buf_final_merged_1_rst), .start(buf_final_merged_1_start), .done(buf_final_merged_1_done), .final_merged_1_update_0_write_wen(buf_final_merged_1_final_merged_1_update_0_write_wen), .final_merged_1_update_0_write_wdata(buf_final_merged_1_final_merged_1_update_0_write_wdata), .final_merged_0_update_0_read_dummy(buf_final_merged_1_final_merged_0_update_0_read_dummy), .final_merged_0_update_0_read_rdata(buf_final_merged_1_final_merged_0_update_0_read_rdata));
  assign buf_final_merged_1_clk = clk;
  assign buf_final_merged_1_rst = rst;
  assign buf_final_merged_1_start = start;
  // Bindings to buf_final_merged_1
    // final_merged_1_final_merged_1_update_0_write_write_122
  assign final_merged_1_final_merged_1_update_0_write_write_122 = buf_final_merged_1_final_merged_1_update_0_write_wdata;
  assign buf_final_merged_1_final_merged_1_update_0_write_wen = stage_172_active;
    // final_merged_1_final_merged_0_update_0_read_read_123
  assign final_merged_1_final_merged_0_update_0_read_read_123 = buf_final_merged_1_final_merged_0_update_0_read_rdata;

  // buf_final_merged_2
  logic [0:0] buf_final_merged_2_clk;
  logic [0:0] buf_final_merged_2_rst;
  logic [0:0] buf_final_merged_2_start;
  logic [0:0] buf_final_merged_2_done;
  logic [31:0] buf_final_merged_2_final_merged_2_update_0_write_wdata;
  logic [0:0] buf_final_merged_2_final_merged_2_update_0_write_wen;
  logic [31:0] buf_final_merged_2_final_merged_1_update_0_read_dummy;
  logic [31:0] buf_final_merged_2_final_merged_1_update_0_read_rdata;
  final_merged_2 buf_final_merged_2(.clk(buf_final_merged_2_clk), .rst(buf_final_merged_2_rst), .start(buf_final_merged_2_start), .done(buf_final_merged_2_done), .final_merged_2_update_0_write_wdata(buf_final_merged_2_final_merged_2_update_0_write_wdata), .final_merged_2_update_0_write_wen(buf_final_merged_2_final_merged_2_update_0_write_wen), .final_merged_1_update_0_read_dummy(buf_final_merged_2_final_merged_1_update_0_read_dummy), .final_merged_1_update_0_read_rdata(buf_final_merged_2_final_merged_1_update_0_read_rdata));
  assign buf_final_merged_2_clk = clk;
  assign buf_final_merged_2_rst = rst;
  assign buf_final_merged_2_start = start;
  // Bindings to buf_final_merged_2
    // final_merged_2_final_merged_1_update_0_read_read_120
  assign final_merged_2_final_merged_1_update_0_read_read_120 = buf_final_merged_2_final_merged_1_update_0_read_rdata;
    // final_merged_2_final_merged_2_update_0_write_write_119
  assign final_merged_2_final_merged_2_update_0_write_write_119 = buf_final_merged_2_final_merged_2_update_0_write_wdata;
  assign buf_final_merged_2_final_merged_2_update_0_write_wen = stage_168_active;

  // buf_fused_level_0
  logic [0:0] buf_fused_level_0_clk;
  logic [0:0] buf_fused_level_0_rst;
  logic [0:0] buf_fused_level_0_start;
  logic [0:0] buf_fused_level_0_done;
  logic [0:0] buf_fused_level_0_fused_level_0_update_0_write_wen;
  logic [31:0] buf_fused_level_0_fused_level_0_update_0_write_wdata;
  logic [31:0] buf_fused_level_0_final_merged_0_update_0_read_dummy;
  logic [31:0] buf_fused_level_0_final_merged_0_update_0_read_rdata;
  fused_level_0 buf_fused_level_0(.clk(buf_fused_level_0_clk), .rst(buf_fused_level_0_rst), .start(buf_fused_level_0_start), .done(buf_fused_level_0_done), .fused_level_0_update_0_write_wen(buf_fused_level_0_fused_level_0_update_0_write_wen), .fused_level_0_update_0_write_wdata(buf_fused_level_0_fused_level_0_update_0_write_wdata), .final_merged_0_update_0_read_dummy(buf_fused_level_0_final_merged_0_update_0_read_dummy), .final_merged_0_update_0_read_rdata(buf_fused_level_0_final_merged_0_update_0_read_rdata));
  assign buf_fused_level_0_clk = clk;
  assign buf_fused_level_0_rst = rst;
  assign buf_fused_level_0_start = start;
  // Bindings to buf_fused_level_0
    // fused_level_0_final_merged_0_update_0_read_read_124
  assign fused_level_0_final_merged_0_update_0_read_read_124 = buf_fused_level_0_final_merged_0_update_0_read_rdata;
    // fused_level_0_fused_level_0_update_0_write_write_81
  assign fused_level_0_fused_level_0_update_0_write_write_81 = buf_fused_level_0_fused_level_0_update_0_write_wdata;
  assign buf_fused_level_0_fused_level_0_update_0_write_wen = stage_117_active;

  // buf_fused_level_1
  logic [0:0] buf_fused_level_1_clk;
  logic [0:0] buf_fused_level_1_rst;
  logic [0:0] buf_fused_level_1_start;
  logic [0:0] buf_fused_level_1_done;
  logic [0:0] buf_fused_level_1_fused_level_1_update_0_write_wen;
  logic [31:0] buf_fused_level_1_fused_level_1_update_0_write_wdata;
  logic [31:0] buf_fused_level_1_final_merged_1_update_0_read_dummy;
  logic [31:0] buf_fused_level_1_final_merged_1_update_0_read_rdata;
  fused_level_1 buf_fused_level_1(.clk(buf_fused_level_1_clk), .rst(buf_fused_level_1_rst), .start(buf_fused_level_1_start), .done(buf_fused_level_1_done), .fused_level_1_update_0_write_wen(buf_fused_level_1_fused_level_1_update_0_write_wen), .fused_level_1_update_0_write_wdata(buf_fused_level_1_fused_level_1_update_0_write_wdata), .final_merged_1_update_0_read_dummy(buf_fused_level_1_final_merged_1_update_0_read_dummy), .final_merged_1_update_0_read_rdata(buf_fused_level_1_final_merged_1_update_0_read_rdata));
  assign buf_fused_level_1_clk = clk;
  assign buf_fused_level_1_rst = rst;
  assign buf_fused_level_1_start = start;
  // Bindings to buf_fused_level_1
    // fused_level_1_final_merged_1_update_0_read_read_121
  assign fused_level_1_final_merged_1_update_0_read_read_121 = buf_fused_level_1_final_merged_1_update_0_read_rdata;
    // fused_level_1_fused_level_1_update_0_write_write_89
  assign fused_level_1_fused_level_1_update_0_write_write_89 = buf_fused_level_1_fused_level_1_update_0_write_wdata;
  assign buf_fused_level_1_fused_level_1_update_0_write_wen = stage_127_active;

  // buf_fused_level_2
  logic [0:0] buf_fused_level_2_clk;
  logic [0:0] buf_fused_level_2_rst;
  logic [0:0] buf_fused_level_2_start;
  logic [0:0] buf_fused_level_2_done;
  logic [0:0] buf_fused_level_2_fused_level_2_update_0_write_wen;
  logic [31:0] buf_fused_level_2_fused_level_2_update_0_write_wdata;
  logic [31:0] buf_fused_level_2_final_merged_2_update_0_read_dummy;
  logic [31:0] buf_fused_level_2_final_merged_2_update_0_read_rdata;
  fused_level_2 buf_fused_level_2(.clk(buf_fused_level_2_clk), .rst(buf_fused_level_2_rst), .start(buf_fused_level_2_start), .done(buf_fused_level_2_done), .fused_level_2_update_0_write_wen(buf_fused_level_2_fused_level_2_update_0_write_wen), .fused_level_2_update_0_write_wdata(buf_fused_level_2_fused_level_2_update_0_write_wdata), .final_merged_2_update_0_read_dummy(buf_fused_level_2_final_merged_2_update_0_read_dummy), .final_merged_2_update_0_read_rdata(buf_fused_level_2_final_merged_2_update_0_read_rdata));
  assign buf_fused_level_2_clk = clk;
  assign buf_fused_level_2_rst = rst;
  assign buf_fused_level_2_start = start;
  // Bindings to buf_fused_level_2
    // fused_level_2_final_merged_2_update_0_read_read_118
  assign fused_level_2_final_merged_2_update_0_read_read_118 = buf_fused_level_2_final_merged_2_update_0_read_rdata;
    // fused_level_2_fused_level_2_update_0_write_write_111
  assign fused_level_2_fused_level_2_update_0_write_write_111 = buf_fused_level_2_fused_level_2_update_0_write_wdata;
  assign buf_fused_level_2_fused_level_2_update_0_write_wen = stage_158_active;

  // buf_fused_level_3
  logic [0:0] buf_fused_level_3_clk;
  logic [0:0] buf_fused_level_3_rst;
  logic [0:0] buf_fused_level_3_start;
  logic [0:0] buf_fused_level_3_done;
  logic [0:0] buf_fused_level_3_fused_level_3_update_0_write_wen;
  logic [31:0] buf_fused_level_3_fused_level_3_update_0_write_wdata;
  logic [31:0] buf_fused_level_3_final_merged_2_update_0_read_dummy;
  logic [31:0] buf_fused_level_3_final_merged_2_update_0_read_rdata;
  fused_level_3 buf_fused_level_3(.clk(buf_fused_level_3_clk), .rst(buf_fused_level_3_rst), .start(buf_fused_level_3_start), .done(buf_fused_level_3_done), .fused_level_3_update_0_write_wen(buf_fused_level_3_fused_level_3_update_0_write_wen), .fused_level_3_update_0_write_wdata(buf_fused_level_3_fused_level_3_update_0_write_wdata), .final_merged_2_update_0_read_dummy(buf_fused_level_3_final_merged_2_update_0_read_dummy), .final_merged_2_update_0_read_rdata(buf_fused_level_3_final_merged_2_update_0_read_rdata));
  assign buf_fused_level_3_clk = clk;
  assign buf_fused_level_3_rst = rst;
  assign buf_fused_level_3_start = start;
  // Bindings to buf_fused_level_3
    // fused_level_3_fused_level_3_update_0_write_write_116
  assign fused_level_3_fused_level_3_update_0_write_write_116 = buf_fused_level_3_fused_level_3_update_0_write_wdata;
  assign buf_fused_level_3_fused_level_3_update_0_write_wen = stage_164_active;
    // fused_level_3_final_merged_2_update_0_read_read_117
  assign fused_level_3_final_merged_2_update_0_read_read_117 = buf_fused_level_3_final_merged_2_update_0_read_rdata;

  // buf_in
  logic [0:0] buf_in_clk;
  logic [0:0] buf_in_rst;
  logic [0:0] buf_in_start;
  logic [0:0] buf_in_done;
  logic [0:0] buf_in_in_update_0_write_wen;
  logic [31:0] buf_in_in_update_0_write_wdata;
  logic [31:0] buf_in_bright_update_0_read_dummy;
  logic [31:0] buf_in_bright_update_0_read_rdata;
  logic [31:0] buf_in_dark_update_0_read_dummy;
  logic [31:0] buf_in_dark_update_0_read_rdata;
  in buf_in(.clk(buf_in_clk), .rst(buf_in_rst), .start(buf_in_start), .done(buf_in_done), .in_update_0_write_wen(buf_in_in_update_0_write_wen), .in_update_0_write_wdata(buf_in_in_update_0_write_wdata), .bright_update_0_read_dummy(buf_in_bright_update_0_read_dummy), .bright_update_0_read_rdata(buf_in_bright_update_0_read_rdata), .dark_update_0_read_dummy(buf_in_dark_update_0_read_dummy), .dark_update_0_read_rdata(buf_in_dark_update_0_read_rdata));
  assign buf_in_clk = clk;
  assign buf_in_rst = rst;
  assign buf_in_start = start;
  // Bindings to buf_in
    // in_in_update_0_write_write_1
  assign in_in_update_0_write_write_1 = buf_in_in_update_0_write_wdata;
  assign buf_in_in_update_0_write_wen = stage_2_active;
    // in_bright_update_0_read_read_2
  assign in_bright_update_0_read_read_2 = buf_in_bright_update_0_read_rdata;
    // in_dark_update_0_read_read_6
  assign in_dark_update_0_read_read_6 = buf_in_dark_update_0_read_rdata;

  // Bindings to buf_in_off_chip
    // in_off_chip_in_update_0_read_read_0
  assign in_off_chip_in_update_0_read_read_0 = buf_in_off_chip_in_update_0_read_rdata;

  // buf_weight_sums
  logic [0:0] buf_weight_sums_clk;
  logic [0:0] buf_weight_sums_rst;
  logic [0:0] buf_weight_sums_start;
  logic [0:0] buf_weight_sums_done;
  logic [0:0] buf_weight_sums_weight_sums_update_0_write_wen;
  logic [31:0] buf_weight_sums_weight_sums_update_0_write_wdata;
  logic [31:0] buf_weight_sums_bright_weights_normed_update_0_read_dummy;
  logic [31:0] buf_weight_sums_bright_weights_normed_update_0_read_rdata;
  logic [31:0] buf_weight_sums_dark_weights_normed_update_0_read_dummy;
  logic [31:0] buf_weight_sums_dark_weights_normed_update_0_read_rdata;
  weight_sums buf_weight_sums(.clk(buf_weight_sums_clk), .rst(buf_weight_sums_rst), .start(buf_weight_sums_start), .done(buf_weight_sums_done), .weight_sums_update_0_write_wen(buf_weight_sums_weight_sums_update_0_write_wen), .weight_sums_update_0_write_wdata(buf_weight_sums_weight_sums_update_0_write_wdata), .bright_weights_normed_update_0_read_dummy(buf_weight_sums_bright_weights_normed_update_0_read_dummy), .bright_weights_normed_update_0_read_rdata(buf_weight_sums_bright_weights_normed_update_0_read_rdata), .dark_weights_normed_update_0_read_dummy(buf_weight_sums_dark_weights_normed_update_0_read_dummy), .dark_weights_normed_update_0_read_rdata(buf_weight_sums_dark_weights_normed_update_0_read_rdata));
  assign buf_weight_sums_clk = clk;
  assign buf_weight_sums_rst = rst;
  assign buf_weight_sums_start = start;
  // Bindings to buf_weight_sums
    // weight_sums_weight_sums_update_0_write_write_24
  assign weight_sums_weight_sums_update_0_write_write_24 = buf_weight_sums_weight_sums_update_0_write_wdata;
  assign buf_weight_sums_weight_sums_update_0_write_wen = stage_36_active;
    // weight_sums_bright_weights_normed_update_0_read_read_49
  assign weight_sums_bright_weights_normed_update_0_read_read_49 = buf_weight_sums_bright_weights_normed_update_0_read_rdata;
    // weight_sums_dark_weights_normed_update_0_read_read_46
  assign weight_sums_dark_weights_normed_update_0_read_read_46 = buf_weight_sums_dark_weights_normed_update_0_read_rdata;

  // Bindings to buf_pyramid_synthetic_exposure_fusion
    // pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127
  assign pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_write_127 = buf_pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_wdata;
  assign buf_pyramid_synthetic_exposure_fusion_pyramid_synthetic_exposure_fusion_update_0_write_wen = stage_179_active;

  // in_update_0_128
  logic [0:0] in_update_0_128_clk;
  logic [0:0] in_update_0_128_rst;
  logic [0:0] in_update_0_128_start;
  logic [0:0] in_update_0_128_done;
  logic [31:0] in_update_0_128_src_in;
  logic [31:0] in_update_0_128_src_out;
  logic [31:0] in_update_0_128_out;
  in_update_0 in_update_0_128(.clk(in_update_0_128_clk), .rst(in_update_0_128_rst), .start(in_update_0_128_start), .done(in_update_0_128_done), .src_in(in_update_0_128_src_in), .src_out(in_update_0_128_src_out), .out(in_update_0_128_out));
  assign in_update_0_128_clk = clk;
  assign in_update_0_128_rst = rst;
  assign in_update_0_128_start = start;
  // Bindings to in_update_0_128
    // in_update_0
  assign in_update_0 = in_update_0_128_out;

  // final_merged_1_update_0_132
  logic [0:0] final_merged_1_update_0_132_clk;
  logic [0:0] final_merged_1_update_0_132_rst;
  logic [0:0] final_merged_1_update_0_132_start;
  logic [0:0] final_merged_1_update_0_132_done;
  logic [31:0] final_merged_1_update_0_132_src_in;
  logic [31:0] final_merged_1_update_0_132_src_out;
  logic [31:0] final_merged_1_update_0_132_out;
  final_merged_1_update_0 final_merged_1_update_0_132(.clk(final_merged_1_update_0_132_clk), .rst(final_merged_1_update_0_132_rst), .start(final_merged_1_update_0_132_start), .done(final_merged_1_update_0_132_done), .src_in(final_merged_1_update_0_132_src_in), .src_out(final_merged_1_update_0_132_src_out), .out(final_merged_1_update_0_132_out));
  assign final_merged_1_update_0_132_clk = clk;
  assign final_merged_1_update_0_132_rst = rst;
  assign final_merged_1_update_0_132_start = start;
  // Bindings to final_merged_1_update_0_132
    // final_merged_1_update_0
  assign final_merged_1_update_0 = final_merged_1_update_0_132_out;

  // dark_weights_normed_gauss_blur_2_update_0_131
  logic [0:0] dark_weights_normed_gauss_blur_2_update_0_131_clk;
  logic [0:0] dark_weights_normed_gauss_blur_2_update_0_131_rst;
  logic [0:0] dark_weights_normed_gauss_blur_2_update_0_131_start;
  logic [0:0] dark_weights_normed_gauss_blur_2_update_0_131_done;
  logic [31:0] dark_weights_normed_gauss_blur_2_update_0_131_src_in;
  logic [31:0] dark_weights_normed_gauss_blur_2_update_0_131_src_out;
  logic [31:0] dark_weights_normed_gauss_blur_2_update_0_131_out;
  dark_weights_normed_gauss_blur_2_update_0 dark_weights_normed_gauss_blur_2_update_0_131(.clk(dark_weights_normed_gauss_blur_2_update_0_131_clk), .rst(dark_weights_normed_gauss_blur_2_update_0_131_rst), .start(dark_weights_normed_gauss_blur_2_update_0_131_start), .done(dark_weights_normed_gauss_blur_2_update_0_131_done), .src_in(dark_weights_normed_gauss_blur_2_update_0_131_src_in), .src_out(dark_weights_normed_gauss_blur_2_update_0_131_src_out), .out(dark_weights_normed_gauss_blur_2_update_0_131_out));
  assign dark_weights_normed_gauss_blur_2_update_0_131_clk = clk;
  assign dark_weights_normed_gauss_blur_2_update_0_131_rst = rst;
  assign dark_weights_normed_gauss_blur_2_update_0_131_start = start;
  // Bindings to dark_weights_normed_gauss_blur_2_update_0_131
    // dark_weights_normed_gauss_blur_2_update_0
  assign dark_weights_normed_gauss_blur_2_update_0 = dark_weights_normed_gauss_blur_2_update_0_131_out;

  // bright_gauss_blur_2_update_0_161
  logic [0:0] bright_gauss_blur_2_update_0_161_clk;
  logic [0:0] bright_gauss_blur_2_update_0_161_rst;
  logic [0:0] bright_gauss_blur_2_update_0_161_start;
  logic [0:0] bright_gauss_blur_2_update_0_161_done;
  logic [31:0] bright_gauss_blur_2_update_0_161_src_in;
  logic [31:0] bright_gauss_blur_2_update_0_161_src_out;
  logic [31:0] bright_gauss_blur_2_update_0_161_out;
  bright_gauss_blur_2_update_0 bright_gauss_blur_2_update_0_161(.clk(bright_gauss_blur_2_update_0_161_clk), .rst(bright_gauss_blur_2_update_0_161_rst), .start(bright_gauss_blur_2_update_0_161_start), .done(bright_gauss_blur_2_update_0_161_done), .src_in(bright_gauss_blur_2_update_0_161_src_in), .src_out(bright_gauss_blur_2_update_0_161_src_out), .out(bright_gauss_blur_2_update_0_161_out));
  assign bright_gauss_blur_2_update_0_161_clk = clk;
  assign bright_gauss_blur_2_update_0_161_rst = rst;
  assign bright_gauss_blur_2_update_0_161_start = start;
  // Bindings to bright_gauss_blur_2_update_0_161
    // bright_gauss_blur_2_update_0
  assign bright_gauss_blur_2_update_0 = bright_gauss_blur_2_update_0_161_out;

  // bright_gauss_blur_3_update_0_164
  logic [0:0] bright_gauss_blur_3_update_0_164_clk;
  logic [0:0] bright_gauss_blur_3_update_0_164_rst;
  logic [0:0] bright_gauss_blur_3_update_0_164_start;
  logic [0:0] bright_gauss_blur_3_update_0_164_done;
  logic [31:0] bright_gauss_blur_3_update_0_164_out;
  logic [31:0] bright_gauss_blur_3_update_0_164_src_in;
  logic [31:0] bright_gauss_blur_3_update_0_164_src_out;
  bright_gauss_blur_3_update_0 bright_gauss_blur_3_update_0_164(.clk(bright_gauss_blur_3_update_0_164_clk), .rst(bright_gauss_blur_3_update_0_164_rst), .start(bright_gauss_blur_3_update_0_164_start), .done(bright_gauss_blur_3_update_0_164_done), .out(bright_gauss_blur_3_update_0_164_out), .src_in(bright_gauss_blur_3_update_0_164_src_in), .src_out(bright_gauss_blur_3_update_0_164_src_out));
  assign bright_gauss_blur_3_update_0_164_clk = clk;
  assign bright_gauss_blur_3_update_0_164_rst = rst;
  assign bright_gauss_blur_3_update_0_164_start = start;
  // Bindings to bright_gauss_blur_3_update_0_164
    // bright_gauss_blur_3_update_0
  assign bright_gauss_blur_3_update_0 = bright_gauss_blur_3_update_0_164_out;

  // bright_laplace_diff_2_update_0_172
  logic [0:0] bright_laplace_diff_2_update_0_172_clk;
  logic [0:0] bright_laplace_diff_2_update_0_172_rst;
  logic [0:0] bright_laplace_diff_2_update_0_172_start;
  logic [0:0] bright_laplace_diff_2_update_0_172_done;
  logic [31:0] bright_laplace_diff_2_update_0_172_src_in;
  logic [31:0] bright_laplace_diff_2_update_0_172_src_out;
  logic [31:0] bright_laplace_diff_2_update_0_172_out;
  bright_laplace_diff_2_update_0 bright_laplace_diff_2_update_0_172(.clk(bright_laplace_diff_2_update_0_172_clk), .rst(bright_laplace_diff_2_update_0_172_rst), .start(bright_laplace_diff_2_update_0_172_start), .done(bright_laplace_diff_2_update_0_172_done), .src_in(bright_laplace_diff_2_update_0_172_src_in), .src_out(bright_laplace_diff_2_update_0_172_src_out), .out(bright_laplace_diff_2_update_0_172_out));
  assign bright_laplace_diff_2_update_0_172_clk = clk;
  assign bright_laplace_diff_2_update_0_172_rst = rst;
  assign bright_laplace_diff_2_update_0_172_start = start;
  // Bindings to bright_laplace_diff_2_update_0_172
    // bright_laplace_diff_2_update_0
  assign bright_laplace_diff_2_update_0 = bright_laplace_diff_2_update_0_172_out;

  // fused_level_0_update_0_171
  logic [0:0] fused_level_0_update_0_171_clk;
  logic [0:0] fused_level_0_update_0_171_rst;
  logic [0:0] fused_level_0_update_0_171_start;
  logic [0:0] fused_level_0_update_0_171_done;
  logic [31:0] fused_level_0_update_0_171_src_in;
  logic [31:0] fused_level_0_update_0_171_src_out;
  logic [31:0] fused_level_0_update_0_171_out;
  fused_level_0_update_0 fused_level_0_update_0_171(.clk(fused_level_0_update_0_171_clk), .rst(fused_level_0_update_0_171_rst), .start(fused_level_0_update_0_171_start), .done(fused_level_0_update_0_171_done), .src_in(fused_level_0_update_0_171_src_in), .src_out(fused_level_0_update_0_171_src_out), .out(fused_level_0_update_0_171_out));
  assign fused_level_0_update_0_171_clk = clk;
  assign fused_level_0_update_0_171_rst = rst;
  assign fused_level_0_update_0_171_start = start;
  // Bindings to fused_level_0_update_0_171
    // fused_level_0_update_0
  assign fused_level_0_update_0 = fused_level_0_update_0_171_out;

  // dark_laplace_diff_2_update_0_176
  logic [0:0] dark_laplace_diff_2_update_0_176_clk;
  logic [0:0] dark_laplace_diff_2_update_0_176_rst;
  logic [0:0] dark_laplace_diff_2_update_0_176_start;
  logic [0:0] dark_laplace_diff_2_update_0_176_done;
  logic [31:0] dark_laplace_diff_2_update_0_176_src_in;
  logic [31:0] dark_laplace_diff_2_update_0_176_src_out;
  logic [31:0] dark_laplace_diff_2_update_0_176_out;
  dark_laplace_diff_2_update_0 dark_laplace_diff_2_update_0_176(.clk(dark_laplace_diff_2_update_0_176_clk), .rst(dark_laplace_diff_2_update_0_176_rst), .start(dark_laplace_diff_2_update_0_176_start), .done(dark_laplace_diff_2_update_0_176_done), .src_in(dark_laplace_diff_2_update_0_176_src_in), .src_out(dark_laplace_diff_2_update_0_176_src_out), .out(dark_laplace_diff_2_update_0_176_out));
  assign dark_laplace_diff_2_update_0_176_clk = clk;
  assign dark_laplace_diff_2_update_0_176_rst = rst;
  assign dark_laplace_diff_2_update_0_176_start = start;
  // Bindings to dark_laplace_diff_2_update_0_176
    // dark_laplace_diff_2_update_0
  assign dark_laplace_diff_2_update_0 = dark_laplace_diff_2_update_0_176_out;

  // dark_laplace_diff_1_update_0_170
  logic [0:0] dark_laplace_diff_1_update_0_170_clk;
  logic [0:0] dark_laplace_diff_1_update_0_170_rst;
  logic [0:0] dark_laplace_diff_1_update_0_170_start;
  logic [0:0] dark_laplace_diff_1_update_0_170_done;
  logic [31:0] dark_laplace_diff_1_update_0_170_out;
  logic [31:0] dark_laplace_diff_1_update_0_170_src_in;
  logic [31:0] dark_laplace_diff_1_update_0_170_src_out;
  dark_laplace_diff_1_update_0 dark_laplace_diff_1_update_0_170(.clk(dark_laplace_diff_1_update_0_170_clk), .rst(dark_laplace_diff_1_update_0_170_rst), .start(dark_laplace_diff_1_update_0_170_start), .done(dark_laplace_diff_1_update_0_170_done), .out(dark_laplace_diff_1_update_0_170_out), .src_in(dark_laplace_diff_1_update_0_170_src_in), .src_out(dark_laplace_diff_1_update_0_170_src_out));
  assign dark_laplace_diff_1_update_0_170_clk = clk;
  assign dark_laplace_diff_1_update_0_170_rst = rst;
  assign dark_laplace_diff_1_update_0_170_start = start;
  // Bindings to dark_laplace_diff_1_update_0_170
    // dark_laplace_diff_1_update_0
  assign dark_laplace_diff_1_update_0 = dark_laplace_diff_1_update_0_170_out;

  // dark_weights_normed_gauss_blur_1_update_0_165
  logic [0:0] dark_weights_normed_gauss_blur_1_update_0_165_clk;
  logic [0:0] dark_weights_normed_gauss_blur_1_update_0_165_rst;
  logic [0:0] dark_weights_normed_gauss_blur_1_update_0_165_start;
  logic [0:0] dark_weights_normed_gauss_blur_1_update_0_165_done;
  logic [31:0] dark_weights_normed_gauss_blur_1_update_0_165_src_in;
  logic [31:0] dark_weights_normed_gauss_blur_1_update_0_165_src_out;
  logic [31:0] dark_weights_normed_gauss_blur_1_update_0_165_out;
  dark_weights_normed_gauss_blur_1_update_0 dark_weights_normed_gauss_blur_1_update_0_165(.clk(dark_weights_normed_gauss_blur_1_update_0_165_clk), .rst(dark_weights_normed_gauss_blur_1_update_0_165_rst), .start(dark_weights_normed_gauss_blur_1_update_0_165_start), .done(dark_weights_normed_gauss_blur_1_update_0_165_done), .src_in(dark_weights_normed_gauss_blur_1_update_0_165_src_in), .src_out(dark_weights_normed_gauss_blur_1_update_0_165_src_out), .out(dark_weights_normed_gauss_blur_1_update_0_165_out));
  assign dark_weights_normed_gauss_blur_1_update_0_165_clk = clk;
  assign dark_weights_normed_gauss_blur_1_update_0_165_rst = rst;
  assign dark_weights_normed_gauss_blur_1_update_0_165_start = start;
  // Bindings to dark_weights_normed_gauss_blur_1_update_0_165
    // dark_weights_normed_gauss_blur_1_update_0
  assign dark_weights_normed_gauss_blur_1_update_0 = dark_weights_normed_gauss_blur_1_update_0_165_out;

  // bright_laplace_diff_1_update_0_168
  logic [0:0] bright_laplace_diff_1_update_0_168_clk;
  logic [0:0] bright_laplace_diff_1_update_0_168_rst;
  logic [0:0] bright_laplace_diff_1_update_0_168_start;
  logic [0:0] bright_laplace_diff_1_update_0_168_done;
  logic [31:0] bright_laplace_diff_1_update_0_168_src_in;
  logic [31:0] bright_laplace_diff_1_update_0_168_src_out;
  logic [31:0] bright_laplace_diff_1_update_0_168_out;
  bright_laplace_diff_1_update_0 bright_laplace_diff_1_update_0_168(.clk(bright_laplace_diff_1_update_0_168_clk), .rst(bright_laplace_diff_1_update_0_168_rst), .start(bright_laplace_diff_1_update_0_168_start), .done(bright_laplace_diff_1_update_0_168_done), .src_in(bright_laplace_diff_1_update_0_168_src_in), .src_out(bright_laplace_diff_1_update_0_168_src_out), .out(bright_laplace_diff_1_update_0_168_out));
  assign bright_laplace_diff_1_update_0_168_clk = clk;
  assign bright_laplace_diff_1_update_0_168_rst = rst;
  assign bright_laplace_diff_1_update_0_168_start = start;
  // Bindings to bright_laplace_diff_1_update_0_168
    // bright_laplace_diff_1_update_0
  assign bright_laplace_diff_1_update_0 = bright_laplace_diff_1_update_0_168_out;

  // dark_weights_normed_gauss_blur_3_update_0_169
  logic [0:0] dark_weights_normed_gauss_blur_3_update_0_169_clk;
  logic [0:0] dark_weights_normed_gauss_blur_3_update_0_169_rst;
  logic [0:0] dark_weights_normed_gauss_blur_3_update_0_169_start;
  logic [0:0] dark_weights_normed_gauss_blur_3_update_0_169_done;
  logic [31:0] dark_weights_normed_gauss_blur_3_update_0_169_src_in;
  logic [31:0] dark_weights_normed_gauss_blur_3_update_0_169_src_out;
  logic [31:0] dark_weights_normed_gauss_blur_3_update_0_169_out;
  dark_weights_normed_gauss_blur_3_update_0 dark_weights_normed_gauss_blur_3_update_0_169(.clk(dark_weights_normed_gauss_blur_3_update_0_169_clk), .rst(dark_weights_normed_gauss_blur_3_update_0_169_rst), .start(dark_weights_normed_gauss_blur_3_update_0_169_start), .done(dark_weights_normed_gauss_blur_3_update_0_169_done), .src_in(dark_weights_normed_gauss_blur_3_update_0_169_src_in), .src_out(dark_weights_normed_gauss_blur_3_update_0_169_src_out), .out(dark_weights_normed_gauss_blur_3_update_0_169_out));
  assign dark_weights_normed_gauss_blur_3_update_0_169_clk = clk;
  assign dark_weights_normed_gauss_blur_3_update_0_169_rst = rst;
  assign dark_weights_normed_gauss_blur_3_update_0_169_start = start;
  // Bindings to dark_weights_normed_gauss_blur_3_update_0_169
    // dark_weights_normed_gauss_blur_3_update_0
  assign dark_weights_normed_gauss_blur_3_update_0 = dark_weights_normed_gauss_blur_3_update_0_169_out;

  // dark_laplace_us_1_update_0_166
  logic [0:0] dark_laplace_us_1_update_0_166_clk;
  logic [0:0] dark_laplace_us_1_update_0_166_rst;
  logic [0:0] dark_laplace_us_1_update_0_166_start;
  logic [0:0] dark_laplace_us_1_update_0_166_done;
  logic [31:0] dark_laplace_us_1_update_0_166_src_in;
  logic [31:0] dark_laplace_us_1_update_0_166_src_out;
  logic [31:0] dark_laplace_us_1_update_0_166_out;
  dark_laplace_us_1_update_0 dark_laplace_us_1_update_0_166(.clk(dark_laplace_us_1_update_0_166_clk), .rst(dark_laplace_us_1_update_0_166_rst), .start(dark_laplace_us_1_update_0_166_start), .done(dark_laplace_us_1_update_0_166_done), .src_in(dark_laplace_us_1_update_0_166_src_in), .src_out(dark_laplace_us_1_update_0_166_src_out), .out(dark_laplace_us_1_update_0_166_out));
  assign dark_laplace_us_1_update_0_166_clk = clk;
  assign dark_laplace_us_1_update_0_166_rst = rst;
  assign dark_laplace_us_1_update_0_166_start = start;
  // Bindings to dark_laplace_us_1_update_0_166
    // dark_laplace_us_1_update_0
  assign dark_laplace_us_1_update_0 = dark_laplace_us_1_update_0_166_out;

  // fused_level_2_update_0_179
  logic [0:0] fused_level_2_update_0_179_clk;
  logic [0:0] fused_level_2_update_0_179_rst;
  logic [0:0] fused_level_2_update_0_179_start;
  logic [0:0] fused_level_2_update_0_179_done;
  logic [31:0] fused_level_2_update_0_179_out;
  logic [31:0] fused_level_2_update_0_179_src_in;
  logic [31:0] fused_level_2_update_0_179_src_out;
  fused_level_2_update_0 fused_level_2_update_0_179(.clk(fused_level_2_update_0_179_clk), .rst(fused_level_2_update_0_179_rst), .start(fused_level_2_update_0_179_start), .done(fused_level_2_update_0_179_done), .out(fused_level_2_update_0_179_out), .src_in(fused_level_2_update_0_179_src_in), .src_out(fused_level_2_update_0_179_src_out));
  assign fused_level_2_update_0_179_clk = clk;
  assign fused_level_2_update_0_179_rst = rst;
  assign fused_level_2_update_0_179_start = start;
  // Bindings to fused_level_2_update_0_179
    // fused_level_2_update_0
  assign fused_level_2_update_0 = fused_level_2_update_0_179_out;

  // bright_weights_normed_gauss_blur_3_update_0_177
  logic [0:0] bright_weights_normed_gauss_blur_3_update_0_177_clk;
  logic [0:0] bright_weights_normed_gauss_blur_3_update_0_177_rst;
  logic [0:0] bright_weights_normed_gauss_blur_3_update_0_177_start;
  logic [0:0] bright_weights_normed_gauss_blur_3_update_0_177_done;
  logic [31:0] bright_weights_normed_gauss_blur_3_update_0_177_src_in;
  logic [31:0] bright_weights_normed_gauss_blur_3_update_0_177_src_out;
  logic [31:0] bright_weights_normed_gauss_blur_3_update_0_177_out;
  bright_weights_normed_gauss_blur_3_update_0 bright_weights_normed_gauss_blur_3_update_0_177(.clk(bright_weights_normed_gauss_blur_3_update_0_177_clk), .rst(bright_weights_normed_gauss_blur_3_update_0_177_rst), .start(bright_weights_normed_gauss_blur_3_update_0_177_start), .done(bright_weights_normed_gauss_blur_3_update_0_177_done), .src_in(bright_weights_normed_gauss_blur_3_update_0_177_src_in), .src_out(bright_weights_normed_gauss_blur_3_update_0_177_src_out), .out(bright_weights_normed_gauss_blur_3_update_0_177_out));
  assign bright_weights_normed_gauss_blur_3_update_0_177_clk = clk;
  assign bright_weights_normed_gauss_blur_3_update_0_177_rst = rst;
  assign bright_weights_normed_gauss_blur_3_update_0_177_start = start;
  // Bindings to bright_weights_normed_gauss_blur_3_update_0_177
    // bright_weights_normed_gauss_blur_3_update_0
  assign bright_weights_normed_gauss_blur_3_update_0 = bright_weights_normed_gauss_blur_3_update_0_177_out;

  // dark_weights_normed_gauss_ds_2_update_0_167
  logic [0:0] dark_weights_normed_gauss_ds_2_update_0_167_clk;
  logic [0:0] dark_weights_normed_gauss_ds_2_update_0_167_rst;
  logic [0:0] dark_weights_normed_gauss_ds_2_update_0_167_start;
  logic [0:0] dark_weights_normed_gauss_ds_2_update_0_167_done;
  logic [31:0] dark_weights_normed_gauss_ds_2_update_0_167_src_in;
  logic [31:0] dark_weights_normed_gauss_ds_2_update_0_167_src_out;
  logic [31:0] dark_weights_normed_gauss_ds_2_update_0_167_out;
  dark_weights_normed_gauss_ds_2_update_0 dark_weights_normed_gauss_ds_2_update_0_167(.clk(dark_weights_normed_gauss_ds_2_update_0_167_clk), .rst(dark_weights_normed_gauss_ds_2_update_0_167_rst), .start(dark_weights_normed_gauss_ds_2_update_0_167_start), .done(dark_weights_normed_gauss_ds_2_update_0_167_done), .src_in(dark_weights_normed_gauss_ds_2_update_0_167_src_in), .src_out(dark_weights_normed_gauss_ds_2_update_0_167_src_out), .out(dark_weights_normed_gauss_ds_2_update_0_167_out));
  assign dark_weights_normed_gauss_ds_2_update_0_167_clk = clk;
  assign dark_weights_normed_gauss_ds_2_update_0_167_rst = rst;
  assign dark_weights_normed_gauss_ds_2_update_0_167_start = start;
  // Bindings to dark_weights_normed_gauss_ds_2_update_0_167
    // dark_weights_normed_gauss_ds_2_update_0
  assign dark_weights_normed_gauss_ds_2_update_0 = dark_weights_normed_gauss_ds_2_update_0_167_out;

  // bright_update_0_133
  logic [0:0] bright_update_0_133_clk;
  logic [0:0] bright_update_0_133_rst;
  logic [0:0] bright_update_0_133_start;
  logic [0:0] bright_update_0_133_done;
  logic [31:0] bright_update_0_133_src_in;
  logic [31:0] bright_update_0_133_src_out;
  logic [31:0] bright_update_0_133_out;
  bright_update_0 bright_update_0_133(.clk(bright_update_0_133_clk), .rst(bright_update_0_133_rst), .start(bright_update_0_133_start), .done(bright_update_0_133_done), .src_in(bright_update_0_133_src_in), .src_out(bright_update_0_133_src_out), .out(bright_update_0_133_out));
  assign bright_update_0_133_clk = clk;
  assign bright_update_0_133_rst = rst;
  assign bright_update_0_133_start = start;
  // Bindings to bright_update_0_133
    // bright_update_0
  assign bright_update_0 = bright_update_0_133_out;

  // bright_weights_update_0_129
  logic [0:0] bright_weights_update_0_129_clk;
  logic [0:0] bright_weights_update_0_129_rst;
  logic [0:0] bright_weights_update_0_129_start;
  logic [0:0] bright_weights_update_0_129_done;
  logic [31:0] bright_weights_update_0_129_src_in;
  logic [31:0] bright_weights_update_0_129_src_out;
  logic [31:0] bright_weights_update_0_129_out;
  bright_weights_update_0 bright_weights_update_0_129(.clk(bright_weights_update_0_129_clk), .rst(bright_weights_update_0_129_rst), .start(bright_weights_update_0_129_start), .done(bright_weights_update_0_129_done), .src_in(bright_weights_update_0_129_src_in), .src_out(bright_weights_update_0_129_src_out), .out(bright_weights_update_0_129_out));
  assign bright_weights_update_0_129_clk = clk;
  assign bright_weights_update_0_129_rst = rst;
  assign bright_weights_update_0_129_start = start;
  // Bindings to bright_weights_update_0_129
    // bright_weights_update_0
  assign bright_weights_update_0 = bright_weights_update_0_129_out;

  // bright_gauss_ds_1_update_0_159
  logic [0:0] bright_gauss_ds_1_update_0_159_clk;
  logic [0:0] bright_gauss_ds_1_update_0_159_rst;
  logic [0:0] bright_gauss_ds_1_update_0_159_start;
  logic [0:0] bright_gauss_ds_1_update_0_159_done;
  logic [31:0] bright_gauss_ds_1_update_0_159_out;
  logic [31:0] bright_gauss_ds_1_update_0_159_src_in;
  logic [31:0] bright_gauss_ds_1_update_0_159_src_out;
  bright_gauss_ds_1_update_0 bright_gauss_ds_1_update_0_159(.clk(bright_gauss_ds_1_update_0_159_clk), .rst(bright_gauss_ds_1_update_0_159_rst), .start(bright_gauss_ds_1_update_0_159_start), .done(bright_gauss_ds_1_update_0_159_done), .out(bright_gauss_ds_1_update_0_159_out), .src_in(bright_gauss_ds_1_update_0_159_src_in), .src_out(bright_gauss_ds_1_update_0_159_src_out));
  assign bright_gauss_ds_1_update_0_159_clk = clk;
  assign bright_gauss_ds_1_update_0_159_rst = rst;
  assign bright_gauss_ds_1_update_0_159_start = start;
  // Bindings to bright_gauss_ds_1_update_0_159
    // bright_gauss_ds_1_update_0
  assign bright_gauss_ds_1_update_0 = bright_gauss_ds_1_update_0_159_out;

  // dark_update_0_134
  logic [0:0] dark_update_0_134_clk;
  logic [0:0] dark_update_0_134_rst;
  logic [0:0] dark_update_0_134_start;
  logic [0:0] dark_update_0_134_done;
  logic [31:0] dark_update_0_134_src_in;
  logic [31:0] dark_update_0_134_src_out;
  logic [31:0] dark_update_0_134_out;
  dark_update_0 dark_update_0_134(.clk(dark_update_0_134_clk), .rst(dark_update_0_134_rst), .start(dark_update_0_134_start), .done(dark_update_0_134_done), .src_in(dark_update_0_134_src_in), .src_out(dark_update_0_134_src_out), .out(dark_update_0_134_out));
  assign dark_update_0_134_clk = clk;
  assign dark_update_0_134_rst = rst;
  assign dark_update_0_134_start = start;
  // Bindings to dark_update_0_134
    // dark_update_0
  assign dark_update_0 = dark_update_0_134_out;

  // dark_gauss_ds_2_update_0_163
  logic [0:0] dark_gauss_ds_2_update_0_163_clk;
  logic [0:0] dark_gauss_ds_2_update_0_163_rst;
  logic [0:0] dark_gauss_ds_2_update_0_163_start;
  logic [0:0] dark_gauss_ds_2_update_0_163_done;
  logic [31:0] dark_gauss_ds_2_update_0_163_src_in;
  logic [31:0] dark_gauss_ds_2_update_0_163_src_out;
  logic [31:0] dark_gauss_ds_2_update_0_163_out;
  dark_gauss_ds_2_update_0 dark_gauss_ds_2_update_0_163(.clk(dark_gauss_ds_2_update_0_163_clk), .rst(dark_gauss_ds_2_update_0_163_rst), .start(dark_gauss_ds_2_update_0_163_start), .done(dark_gauss_ds_2_update_0_163_done), .src_in(dark_gauss_ds_2_update_0_163_src_in), .src_out(dark_gauss_ds_2_update_0_163_src_out), .out(dark_gauss_ds_2_update_0_163_out));
  assign dark_gauss_ds_2_update_0_163_clk = clk;
  assign dark_gauss_ds_2_update_0_163_rst = rst;
  assign dark_gauss_ds_2_update_0_163_start = start;
  // Bindings to dark_gauss_ds_2_update_0_163
    // dark_gauss_ds_2_update_0
  assign dark_gauss_ds_2_update_0 = dark_gauss_ds_2_update_0_163_out;

  // dark_weights_update_0_130
  logic [0:0] dark_weights_update_0_130_clk;
  logic [0:0] dark_weights_update_0_130_rst;
  logic [0:0] dark_weights_update_0_130_start;
  logic [0:0] dark_weights_update_0_130_done;
  logic [31:0] dark_weights_update_0_130_src_in;
  logic [31:0] dark_weights_update_0_130_src_out;
  logic [31:0] dark_weights_update_0_130_out;
  dark_weights_update_0 dark_weights_update_0_130(.clk(dark_weights_update_0_130_clk), .rst(dark_weights_update_0_130_rst), .start(dark_weights_update_0_130_start), .done(dark_weights_update_0_130_done), .src_in(dark_weights_update_0_130_src_in), .src_out(dark_weights_update_0_130_src_out), .out(dark_weights_update_0_130_out));
  assign dark_weights_update_0_130_clk = clk;
  assign dark_weights_update_0_130_rst = rst;
  assign dark_weights_update_0_130_start = start;
  // Bindings to dark_weights_update_0_130
    // dark_weights_update_0
  assign dark_weights_update_0 = dark_weights_update_0_130_out;

  // dark_gauss_blur_3_update_0_151
  logic [0:0] dark_gauss_blur_3_update_0_151_clk;
  logic [0:0] dark_gauss_blur_3_update_0_151_rst;
  logic [0:0] dark_gauss_blur_3_update_0_151_start;
  logic [0:0] dark_gauss_blur_3_update_0_151_done;
  logic [31:0] dark_gauss_blur_3_update_0_151_src_in;
  logic [31:0] dark_gauss_blur_3_update_0_151_src_out;
  logic [31:0] dark_gauss_blur_3_update_0_151_out;
  dark_gauss_blur_3_update_0 dark_gauss_blur_3_update_0_151(.clk(dark_gauss_blur_3_update_0_151_clk), .rst(dark_gauss_blur_3_update_0_151_rst), .start(dark_gauss_blur_3_update_0_151_start), .done(dark_gauss_blur_3_update_0_151_done), .src_in(dark_gauss_blur_3_update_0_151_src_in), .src_out(dark_gauss_blur_3_update_0_151_src_out), .out(dark_gauss_blur_3_update_0_151_out));
  assign dark_gauss_blur_3_update_0_151_clk = clk;
  assign dark_gauss_blur_3_update_0_151_rst = rst;
  assign dark_gauss_blur_3_update_0_151_start = start;
  // Bindings to dark_gauss_blur_3_update_0_151
    // dark_gauss_blur_3_update_0
  assign dark_gauss_blur_3_update_0 = dark_gauss_blur_3_update_0_151_out;

  // bright_gauss_ds_3_update_0_147
  logic [0:0] bright_gauss_ds_3_update_0_147_clk;
  logic [0:0] bright_gauss_ds_3_update_0_147_rst;
  logic [0:0] bright_gauss_ds_3_update_0_147_start;
  logic [0:0] bright_gauss_ds_3_update_0_147_done;
  logic [31:0] bright_gauss_ds_3_update_0_147_src_in;
  logic [31:0] bright_gauss_ds_3_update_0_147_src_out;
  logic [31:0] bright_gauss_ds_3_update_0_147_out;
  bright_gauss_ds_3_update_0 bright_gauss_ds_3_update_0_147(.clk(bright_gauss_ds_3_update_0_147_clk), .rst(bright_gauss_ds_3_update_0_147_rst), .start(bright_gauss_ds_3_update_0_147_start), .done(bright_gauss_ds_3_update_0_147_done), .src_in(bright_gauss_ds_3_update_0_147_src_in), .src_out(bright_gauss_ds_3_update_0_147_src_out), .out(bright_gauss_ds_3_update_0_147_out));
  assign bright_gauss_ds_3_update_0_147_clk = clk;
  assign bright_gauss_ds_3_update_0_147_rst = rst;
  assign bright_gauss_ds_3_update_0_147_start = start;
  // Bindings to bright_gauss_ds_3_update_0_147
    // bright_gauss_ds_3_update_0
  assign bright_gauss_ds_3_update_0 = bright_gauss_ds_3_update_0_147_out;

  // bright_weights_normed_gauss_ds_3_update_0_178
  logic [0:0] bright_weights_normed_gauss_ds_3_update_0_178_clk;
  logic [0:0] bright_weights_normed_gauss_ds_3_update_0_178_rst;
  logic [0:0] bright_weights_normed_gauss_ds_3_update_0_178_start;
  logic [0:0] bright_weights_normed_gauss_ds_3_update_0_178_done;
  logic [31:0] bright_weights_normed_gauss_ds_3_update_0_178_src_in;
  logic [31:0] bright_weights_normed_gauss_ds_3_update_0_178_src_out;
  logic [31:0] bright_weights_normed_gauss_ds_3_update_0_178_out;
  bright_weights_normed_gauss_ds_3_update_0 bright_weights_normed_gauss_ds_3_update_0_178(.clk(bright_weights_normed_gauss_ds_3_update_0_178_clk), .rst(bright_weights_normed_gauss_ds_3_update_0_178_rst), .start(bright_weights_normed_gauss_ds_3_update_0_178_start), .done(bright_weights_normed_gauss_ds_3_update_0_178_done), .src_in(bright_weights_normed_gauss_ds_3_update_0_178_src_in), .src_out(bright_weights_normed_gauss_ds_3_update_0_178_src_out), .out(bright_weights_normed_gauss_ds_3_update_0_178_out));
  assign bright_weights_normed_gauss_ds_3_update_0_178_clk = clk;
  assign bright_weights_normed_gauss_ds_3_update_0_178_rst = rst;
  assign bright_weights_normed_gauss_ds_3_update_0_178_start = start;
  // Bindings to bright_weights_normed_gauss_ds_3_update_0_178
    // bright_weights_normed_gauss_ds_3_update_0
  assign bright_weights_normed_gauss_ds_3_update_0 = bright_weights_normed_gauss_ds_3_update_0_178_out;

  // dark_gauss_blur_2_update_0_158
  logic [0:0] dark_gauss_blur_2_update_0_158_clk;
  logic [0:0] dark_gauss_blur_2_update_0_158_rst;
  logic [0:0] dark_gauss_blur_2_update_0_158_start;
  logic [0:0] dark_gauss_blur_2_update_0_158_done;
  logic [31:0] dark_gauss_blur_2_update_0_158_src_in;
  logic [31:0] dark_gauss_blur_2_update_0_158_src_out;
  logic [31:0] dark_gauss_blur_2_update_0_158_out;
  dark_gauss_blur_2_update_0 dark_gauss_blur_2_update_0_158(.clk(dark_gauss_blur_2_update_0_158_clk), .rst(dark_gauss_blur_2_update_0_158_rst), .start(dark_gauss_blur_2_update_0_158_start), .done(dark_gauss_blur_2_update_0_158_done), .src_in(dark_gauss_blur_2_update_0_158_src_in), .src_out(dark_gauss_blur_2_update_0_158_src_out), .out(dark_gauss_blur_2_update_0_158_out));
  assign dark_gauss_blur_2_update_0_158_clk = clk;
  assign dark_gauss_blur_2_update_0_158_rst = rst;
  assign dark_gauss_blur_2_update_0_158_start = start;
  // Bindings to dark_gauss_blur_2_update_0_158
    // dark_gauss_blur_2_update_0
  assign dark_gauss_blur_2_update_0 = dark_gauss_blur_2_update_0_158_out;

  // dark_gauss_ds_1_update_0_157
  logic [0:0] dark_gauss_ds_1_update_0_157_clk;
  logic [0:0] dark_gauss_ds_1_update_0_157_rst;
  logic [0:0] dark_gauss_ds_1_update_0_157_start;
  logic [0:0] dark_gauss_ds_1_update_0_157_done;
  logic [31:0] dark_gauss_ds_1_update_0_157_src_in;
  logic [31:0] dark_gauss_ds_1_update_0_157_src_out;
  logic [31:0] dark_gauss_ds_1_update_0_157_out;
  dark_gauss_ds_1_update_0 dark_gauss_ds_1_update_0_157(.clk(dark_gauss_ds_1_update_0_157_clk), .rst(dark_gauss_ds_1_update_0_157_rst), .start(dark_gauss_ds_1_update_0_157_start), .done(dark_gauss_ds_1_update_0_157_done), .src_in(dark_gauss_ds_1_update_0_157_src_in), .src_out(dark_gauss_ds_1_update_0_157_src_out), .out(dark_gauss_ds_1_update_0_157_out));
  assign dark_gauss_ds_1_update_0_157_clk = clk;
  assign dark_gauss_ds_1_update_0_157_rst = rst;
  assign dark_gauss_ds_1_update_0_157_start = start;
  // Bindings to dark_gauss_ds_1_update_0_157
    // dark_gauss_ds_1_update_0
  assign dark_gauss_ds_1_update_0 = dark_gauss_ds_1_update_0_157_out;

  // dark_laplace_us_2_update_0_155
  logic [0:0] dark_laplace_us_2_update_0_155_clk;
  logic [0:0] dark_laplace_us_2_update_0_155_rst;
  logic [0:0] dark_laplace_us_2_update_0_155_start;
  logic [0:0] dark_laplace_us_2_update_0_155_done;
  logic [31:0] dark_laplace_us_2_update_0_155_src_in;
  logic [31:0] dark_laplace_us_2_update_0_155_src_out;
  logic [31:0] dark_laplace_us_2_update_0_155_out;
  dark_laplace_us_2_update_0 dark_laplace_us_2_update_0_155(.clk(dark_laplace_us_2_update_0_155_clk), .rst(dark_laplace_us_2_update_0_155_rst), .start(dark_laplace_us_2_update_0_155_start), .done(dark_laplace_us_2_update_0_155_done), .src_in(dark_laplace_us_2_update_0_155_src_in), .src_out(dark_laplace_us_2_update_0_155_src_out), .out(dark_laplace_us_2_update_0_155_out));
  assign dark_laplace_us_2_update_0_155_clk = clk;
  assign dark_laplace_us_2_update_0_155_rst = rst;
  assign dark_laplace_us_2_update_0_155_start = start;
  // Bindings to dark_laplace_us_2_update_0_155
    // dark_laplace_us_2_update_0
  assign dark_laplace_us_2_update_0 = dark_laplace_us_2_update_0_155_out;

  // fused_level_1_update_0_153
  logic [0:0] fused_level_1_update_0_153_clk;
  logic [0:0] fused_level_1_update_0_153_rst;
  logic [0:0] fused_level_1_update_0_153_start;
  logic [0:0] fused_level_1_update_0_153_done;
  logic [31:0] fused_level_1_update_0_153_src_in;
  logic [31:0] fused_level_1_update_0_153_src_out;
  logic [31:0] fused_level_1_update_0_153_out;
  fused_level_1_update_0 fused_level_1_update_0_153(.clk(fused_level_1_update_0_153_clk), .rst(fused_level_1_update_0_153_rst), .start(fused_level_1_update_0_153_start), .done(fused_level_1_update_0_153_done), .src_in(fused_level_1_update_0_153_src_in), .src_out(fused_level_1_update_0_153_src_out), .out(fused_level_1_update_0_153_out));
  assign fused_level_1_update_0_153_clk = clk;
  assign fused_level_1_update_0_153_rst = rst;
  assign fused_level_1_update_0_153_start = start;
  // Bindings to fused_level_1_update_0_153
    // fused_level_1_update_0
  assign fused_level_1_update_0 = fused_level_1_update_0_153_out;

  // bright_weights_normed_gauss_ds_1_update_0_152
  logic [0:0] bright_weights_normed_gauss_ds_1_update_0_152_clk;
  logic [0:0] bright_weights_normed_gauss_ds_1_update_0_152_rst;
  logic [0:0] bright_weights_normed_gauss_ds_1_update_0_152_start;
  logic [0:0] bright_weights_normed_gauss_ds_1_update_0_152_done;
  logic [31:0] bright_weights_normed_gauss_ds_1_update_0_152_src_in;
  logic [31:0] bright_weights_normed_gauss_ds_1_update_0_152_src_out;
  logic [31:0] bright_weights_normed_gauss_ds_1_update_0_152_out;
  bright_weights_normed_gauss_ds_1_update_0 bright_weights_normed_gauss_ds_1_update_0_152(.clk(bright_weights_normed_gauss_ds_1_update_0_152_clk), .rst(bright_weights_normed_gauss_ds_1_update_0_152_rst), .start(bright_weights_normed_gauss_ds_1_update_0_152_start), .done(bright_weights_normed_gauss_ds_1_update_0_152_done), .src_in(bright_weights_normed_gauss_ds_1_update_0_152_src_in), .src_out(bright_weights_normed_gauss_ds_1_update_0_152_src_out), .out(bright_weights_normed_gauss_ds_1_update_0_152_out));
  assign bright_weights_normed_gauss_ds_1_update_0_152_clk = clk;
  assign bright_weights_normed_gauss_ds_1_update_0_152_rst = rst;
  assign bright_weights_normed_gauss_ds_1_update_0_152_start = start;
  // Bindings to bright_weights_normed_gauss_ds_1_update_0_152
    // bright_weights_normed_gauss_ds_1_update_0
  assign bright_weights_normed_gauss_ds_1_update_0 = bright_weights_normed_gauss_ds_1_update_0_152_out;

  // dark_gauss_blur_1_update_0_135
  logic [0:0] dark_gauss_blur_1_update_0_135_clk;
  logic [0:0] dark_gauss_blur_1_update_0_135_rst;
  logic [0:0] dark_gauss_blur_1_update_0_135_start;
  logic [0:0] dark_gauss_blur_1_update_0_135_done;
  logic [31:0] dark_gauss_blur_1_update_0_135_src_in;
  logic [31:0] dark_gauss_blur_1_update_0_135_src_out;
  logic [31:0] dark_gauss_blur_1_update_0_135_out;
  dark_gauss_blur_1_update_0 dark_gauss_blur_1_update_0_135(.clk(dark_gauss_blur_1_update_0_135_clk), .rst(dark_gauss_blur_1_update_0_135_rst), .start(dark_gauss_blur_1_update_0_135_start), .done(dark_gauss_blur_1_update_0_135_done), .src_in(dark_gauss_blur_1_update_0_135_src_in), .src_out(dark_gauss_blur_1_update_0_135_src_out), .out(dark_gauss_blur_1_update_0_135_out));
  assign dark_gauss_blur_1_update_0_135_clk = clk;
  assign dark_gauss_blur_1_update_0_135_rst = rst;
  assign dark_gauss_blur_1_update_0_135_start = start;
  // Bindings to dark_gauss_blur_1_update_0_135
    // dark_gauss_blur_1_update_0
  assign dark_gauss_blur_1_update_0 = dark_gauss_blur_1_update_0_135_out;

  // bright_weights_normed_update_0_149
  logic [0:0] bright_weights_normed_update_0_149_clk;
  logic [0:0] bright_weights_normed_update_0_149_rst;
  logic [0:0] bright_weights_normed_update_0_149_start;
  logic [0:0] bright_weights_normed_update_0_149_done;
  logic [31:0] bright_weights_normed_update_0_149_src_in;
  logic [31:0] bright_weights_normed_update_0_149_src_out;
  logic [31:0] bright_weights_normed_update_0_149_out;
  bright_weights_normed_update_0 bright_weights_normed_update_0_149(.clk(bright_weights_normed_update_0_149_clk), .rst(bright_weights_normed_update_0_149_rst), .start(bright_weights_normed_update_0_149_start), .done(bright_weights_normed_update_0_149_done), .src_in(bright_weights_normed_update_0_149_src_in), .src_out(bright_weights_normed_update_0_149_src_out), .out(bright_weights_normed_update_0_149_out));
  assign bright_weights_normed_update_0_149_clk = clk;
  assign bright_weights_normed_update_0_149_rst = rst;
  assign bright_weights_normed_update_0_149_start = start;
  // Bindings to bright_weights_normed_update_0_149
    // bright_weights_normed_update_0
  assign bright_weights_normed_update_0 = bright_weights_normed_update_0_149_out;

  // bright_gauss_blur_1_update_0_136
  logic [0:0] bright_gauss_blur_1_update_0_136_clk;
  logic [0:0] bright_gauss_blur_1_update_0_136_rst;
  logic [0:0] bright_gauss_blur_1_update_0_136_start;
  logic [0:0] bright_gauss_blur_1_update_0_136_done;
  logic [31:0] bright_gauss_blur_1_update_0_136_src_in;
  logic [31:0] bright_gauss_blur_1_update_0_136_src_out;
  logic [31:0] bright_gauss_blur_1_update_0_136_out;
  bright_gauss_blur_1_update_0 bright_gauss_blur_1_update_0_136(.clk(bright_gauss_blur_1_update_0_136_clk), .rst(bright_gauss_blur_1_update_0_136_rst), .start(bright_gauss_blur_1_update_0_136_start), .done(bright_gauss_blur_1_update_0_136_done), .src_in(bright_gauss_blur_1_update_0_136_src_in), .src_out(bright_gauss_blur_1_update_0_136_src_out), .out(bright_gauss_blur_1_update_0_136_out));
  assign bright_gauss_blur_1_update_0_136_clk = clk;
  assign bright_gauss_blur_1_update_0_136_rst = rst;
  assign bright_gauss_blur_1_update_0_136_start = start;
  // Bindings to bright_gauss_blur_1_update_0_136
    // bright_gauss_blur_1_update_0
  assign bright_gauss_blur_1_update_0 = bright_gauss_blur_1_update_0_136_out;

  // bright_gauss_ds_2_update_0_146
  logic [0:0] bright_gauss_ds_2_update_0_146_clk;
  logic [0:0] bright_gauss_ds_2_update_0_146_rst;
  logic [0:0] bright_gauss_ds_2_update_0_146_start;
  logic [0:0] bright_gauss_ds_2_update_0_146_done;
  logic [31:0] bright_gauss_ds_2_update_0_146_src_in;
  logic [31:0] bright_gauss_ds_2_update_0_146_src_out;
  logic [31:0] bright_gauss_ds_2_update_0_146_out;
  bright_gauss_ds_2_update_0 bright_gauss_ds_2_update_0_146(.clk(bright_gauss_ds_2_update_0_146_clk), .rst(bright_gauss_ds_2_update_0_146_rst), .start(bright_gauss_ds_2_update_0_146_start), .done(bright_gauss_ds_2_update_0_146_done), .src_in(bright_gauss_ds_2_update_0_146_src_in), .src_out(bright_gauss_ds_2_update_0_146_src_out), .out(bright_gauss_ds_2_update_0_146_out));
  assign bright_gauss_ds_2_update_0_146_clk = clk;
  assign bright_gauss_ds_2_update_0_146_rst = rst;
  assign bright_gauss_ds_2_update_0_146_start = start;
  // Bindings to bright_gauss_ds_2_update_0_146
    // bright_gauss_ds_2_update_0
  assign bright_gauss_ds_2_update_0 = bright_gauss_ds_2_update_0_146_out;

  // dark_weights_normed_gauss_ds_3_update_0_154
  logic [0:0] dark_weights_normed_gauss_ds_3_update_0_154_clk;
  logic [0:0] dark_weights_normed_gauss_ds_3_update_0_154_rst;
  logic [0:0] dark_weights_normed_gauss_ds_3_update_0_154_start;
  logic [0:0] dark_weights_normed_gauss_ds_3_update_0_154_done;
  logic [31:0] dark_weights_normed_gauss_ds_3_update_0_154_src_in;
  logic [31:0] dark_weights_normed_gauss_ds_3_update_0_154_src_out;
  logic [31:0] dark_weights_normed_gauss_ds_3_update_0_154_out;
  dark_weights_normed_gauss_ds_3_update_0 dark_weights_normed_gauss_ds_3_update_0_154(.clk(dark_weights_normed_gauss_ds_3_update_0_154_clk), .rst(dark_weights_normed_gauss_ds_3_update_0_154_rst), .start(dark_weights_normed_gauss_ds_3_update_0_154_start), .done(dark_weights_normed_gauss_ds_3_update_0_154_done), .src_in(dark_weights_normed_gauss_ds_3_update_0_154_src_in), .src_out(dark_weights_normed_gauss_ds_3_update_0_154_src_out), .out(dark_weights_normed_gauss_ds_3_update_0_154_out));
  assign dark_weights_normed_gauss_ds_3_update_0_154_clk = clk;
  assign dark_weights_normed_gauss_ds_3_update_0_154_rst = rst;
  assign dark_weights_normed_gauss_ds_3_update_0_154_start = start;
  // Bindings to dark_weights_normed_gauss_ds_3_update_0_154
    // dark_weights_normed_gauss_ds_3_update_0
  assign dark_weights_normed_gauss_ds_3_update_0 = dark_weights_normed_gauss_ds_3_update_0_154_out;

  // bright_laplace_us_0_update_0_162
  logic [0:0] bright_laplace_us_0_update_0_162_clk;
  logic [0:0] bright_laplace_us_0_update_0_162_rst;
  logic [0:0] bright_laplace_us_0_update_0_162_start;
  logic [0:0] bright_laplace_us_0_update_0_162_done;
  logic [31:0] bright_laplace_us_0_update_0_162_src_in;
  logic [31:0] bright_laplace_us_0_update_0_162_src_out;
  logic [31:0] bright_laplace_us_0_update_0_162_out;
  bright_laplace_us_0_update_0 bright_laplace_us_0_update_0_162(.clk(bright_laplace_us_0_update_0_162_clk), .rst(bright_laplace_us_0_update_0_162_rst), .start(bright_laplace_us_0_update_0_162_start), .done(bright_laplace_us_0_update_0_162_done), .src_in(bright_laplace_us_0_update_0_162_src_in), .src_out(bright_laplace_us_0_update_0_162_src_out), .out(bright_laplace_us_0_update_0_162_out));
  assign bright_laplace_us_0_update_0_162_clk = clk;
  assign bright_laplace_us_0_update_0_162_rst = rst;
  assign bright_laplace_us_0_update_0_162_start = start;
  // Bindings to bright_laplace_us_0_update_0_162
    // bright_laplace_us_0_update_0
  assign bright_laplace_us_0_update_0 = bright_laplace_us_0_update_0_162_out;

  // pyramid_synthetic_exposure_fusion_update_0_156
  logic [0:0] pyramid_synthetic_exposure_fusion_update_0_156_clk;
  logic [0:0] pyramid_synthetic_exposure_fusion_update_0_156_rst;
  logic [0:0] pyramid_synthetic_exposure_fusion_update_0_156_start;
  logic [0:0] pyramid_synthetic_exposure_fusion_update_0_156_done;
  logic [31:0] pyramid_synthetic_exposure_fusion_update_0_156_src_in;
  logic [31:0] pyramid_synthetic_exposure_fusion_update_0_156_src_out;
  logic [31:0] pyramid_synthetic_exposure_fusion_update_0_156_out;
  pyramid_synthetic_exposure_fusion_update_0 pyramid_synthetic_exposure_fusion_update_0_156(.clk(pyramid_synthetic_exposure_fusion_update_0_156_clk), .rst(pyramid_synthetic_exposure_fusion_update_0_156_rst), .start(pyramid_synthetic_exposure_fusion_update_0_156_start), .done(pyramid_synthetic_exposure_fusion_update_0_156_done), .src_in(pyramid_synthetic_exposure_fusion_update_0_156_src_in), .src_out(pyramid_synthetic_exposure_fusion_update_0_156_src_out), .out(pyramid_synthetic_exposure_fusion_update_0_156_out));
  assign pyramid_synthetic_exposure_fusion_update_0_156_clk = clk;
  assign pyramid_synthetic_exposure_fusion_update_0_156_rst = rst;
  assign pyramid_synthetic_exposure_fusion_update_0_156_start = start;
  // Bindings to pyramid_synthetic_exposure_fusion_update_0_156
    // pyramid_synthetic_exposure_fusion_update_0
  assign pyramid_synthetic_exposure_fusion_update_0 = pyramid_synthetic_exposure_fusion_update_0_156_out;

  // dark_weights_normed_update_0_160
  logic [0:0] dark_weights_normed_update_0_160_clk;
  logic [0:0] dark_weights_normed_update_0_160_rst;
  logic [0:0] dark_weights_normed_update_0_160_start;
  logic [0:0] dark_weights_normed_update_0_160_done;
  logic [31:0] dark_weights_normed_update_0_160_out;
  logic [31:0] dark_weights_normed_update_0_160_src_in;
  logic [31:0] dark_weights_normed_update_0_160_src_out;
  dark_weights_normed_update_0 dark_weights_normed_update_0_160(.clk(dark_weights_normed_update_0_160_clk), .rst(dark_weights_normed_update_0_160_rst), .start(dark_weights_normed_update_0_160_start), .done(dark_weights_normed_update_0_160_done), .out(dark_weights_normed_update_0_160_out), .src_in(dark_weights_normed_update_0_160_src_in), .src_out(dark_weights_normed_update_0_160_src_out));
  assign dark_weights_normed_update_0_160_clk = clk;
  assign dark_weights_normed_update_0_160_rst = rst;
  assign dark_weights_normed_update_0_160_start = start;
  // Bindings to dark_weights_normed_update_0_160
    // dark_weights_normed_update_0
  assign dark_weights_normed_update_0 = dark_weights_normed_update_0_160_out;


endmodule
