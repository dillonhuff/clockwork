// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U167 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U169 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U156 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U157 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U158 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U160 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U331 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U332 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U327 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U328 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U329 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U330 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U27 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U28 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U23 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U24 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U25 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U26 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U295 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U296 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U291 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U292 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U293 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U294 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U218 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U220 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U206 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U207 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U208 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U210 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U71 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U73 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U59 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U60 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U61 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U63 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U123 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U125 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U111 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U112 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U113 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U115 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U249 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U250 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U245 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U246 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U247 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U248 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U272 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U273 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U268 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U269 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U270 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U271 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module hcompute_hw_output_stencil (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
assign out_hw_output_stencil = in0_conv_stencil[0];
endmodule

module hcompute_hw_kernel_global_wrapper_stencil (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
assign out_hw_kernel_global_wrapper_stencil = in0_hw_kernel_stencil[0];
endmodule

module hcompute_hw_input_global_wrapper_stencil (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
assign out_hw_input_global_wrapper_stencil = in0_hw_input_stencil[0];
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(clk),
    .in(in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire [15:0] enMux_out;
assign enMux_out = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(clk),
    .in(enMux_out),
    .out(out)
);
endmodule

module hcompute_conv_stencil_2 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_1 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_5 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_4 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_3 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U75 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U76_out;
wire [15:0] _U77_out;
wire [15:0] _U78_out;
wire [15:0] _U79_out;
wire [15:0] _U80_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U76 (
    .in(in[0]),
    .clk(clk),
    .out(_U76_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(in[1]),
    .clk(clk),
    .out(_U77_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U78 (
    .in(in[2]),
    .clk(clk),
    .out(_U78_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(in[3]),
    .clk(clk),
    .out(_U79_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(in[4]),
    .clk(clk),
    .out(_U80_out)
);
assign out[4] = _U80_out;
assign out[3] = _U79_out;
assign out[2] = _U78_out;
assign out[1] = _U77_out;
assign out[0] = _U76_out;
endmodule

module array_delay_U65 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U66_out;
wire [15:0] _U67_out;
wire [15:0] _U68_out;
wire [15:0] _U69_out;
wire [15:0] _U70_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(in[0]),
    .clk(clk),
    .out(_U66_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U67 (
    .in(in[1]),
    .clk(clk),
    .out(_U67_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U68 (
    .in(in[2]),
    .clk(clk),
    .out(_U68_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(in[3]),
    .clk(clk),
    .out(_U69_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U70 (
    .in(in[4]),
    .clk(clk),
    .out(_U70_out)
);
assign out[4] = _U70_out;
assign out[3] = _U69_out;
assign out[2] = _U68_out;
assign out[1] = _U67_out;
assign out[0] = _U66_out;
endmodule

module array_delay_U222 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U223_out;
wire [15:0] _U224_out;
wire [15:0] _U225_out;
wire [15:0] _U226_out;
wire [15:0] _U227_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(in[0]),
    .clk(clk),
    .out(_U223_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(in[1]),
    .clk(clk),
    .out(_U224_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(in[2]),
    .clk(clk),
    .out(_U225_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(in[3]),
    .clk(clk),
    .out(_U226_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(in[4]),
    .clk(clk),
    .out(_U227_out)
);
assign out[4] = _U227_out;
assign out[3] = _U226_out;
assign out[2] = _U225_out;
assign out[1] = _U224_out;
assign out[0] = _U223_out;
endmodule

module array_delay_U212 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U213_out;
wire [15:0] _U214_out;
wire [15:0] _U215_out;
wire [15:0] _U216_out;
wire [15:0] _U217_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(in[0]),
    .clk(clk),
    .out(_U213_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(in[1]),
    .clk(clk),
    .out(_U214_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(in[2]),
    .clk(clk),
    .out(_U215_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(in[3]),
    .clk(clk),
    .out(_U216_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(in[4]),
    .clk(clk),
    .out(_U217_out)
);
assign out[4] = _U217_out;
assign out[3] = _U216_out;
assign out[2] = _U215_out;
assign out[1] = _U214_out;
assign out[0] = _U213_out;
endmodule

module array_delay_U171 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U172_out;
wire [15:0] _U173_out;
wire [15:0] _U174_out;
wire [15:0] _U175_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(in[0]),
    .clk(clk),
    .out(_U172_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U173 (
    .in(in[1]),
    .clk(clk),
    .out(_U173_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(in[2]),
    .clk(clk),
    .out(_U174_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(in[3]),
    .clk(clk),
    .out(_U175_out)
);
assign out[3] = _U175_out;
assign out[2] = _U174_out;
assign out[1] = _U173_out;
assign out[0] = _U172_out;
endmodule

module array_delay_U162 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U163_out;
wire [15:0] _U164_out;
wire [15:0] _U165_out;
wire [15:0] _U166_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(in[0]),
    .clk(clk),
    .out(_U163_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(in[1]),
    .clk(clk),
    .out(_U164_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(in[2]),
    .clk(clk),
    .out(_U165_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(in[3]),
    .clk(clk),
    .out(_U166_out)
);
assign out[3] = _U166_out;
assign out[2] = _U165_out;
assign out[1] = _U164_out;
assign out[0] = _U163_out;
endmodule

module array_delay_U127 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U128_out;
wire [15:0] _U129_out;
wire [15:0] _U130_out;
wire [15:0] _U131_out;
wire [15:0] _U132_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(in[0]),
    .clk(clk),
    .out(_U128_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(in[1]),
    .clk(clk),
    .out(_U129_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(in[2]),
    .clk(clk),
    .out(_U130_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U131 (
    .in(in[3]),
    .clk(clk),
    .out(_U131_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(in[4]),
    .clk(clk),
    .out(_U132_out)
);
assign out[4] = _U132_out;
assign out[3] = _U131_out;
assign out[2] = _U130_out;
assign out[1] = _U129_out;
assign out[0] = _U128_out;
endmodule

module array_delay_U117 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U118_out;
wire [15:0] _U119_out;
wire [15:0] _U120_out;
wire [15:0] _U121_out;
wire [15:0] _U122_out;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U118 (
    .in(in[0]),
    .clk(clk),
    .out(_U118_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U119 (
    .in(in[1]),
    .clk(clk),
    .out(_U119_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(in[2]),
    .clk(clk),
    .out(_U120_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U121 (
    .in(in[3]),
    .clk(clk),
    .out(_U121_out)
);
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U122 (
    .in(in[4]),
    .clk(clk),
    .out(_U122_out)
);
assign out[4] = _U122_out;
assign out[3] = _U121_out;
assign out[2] = _U120_out;
assign out[1] = _U119_out;
assign out[0] = _U118_out;
endmodule

module aff__U82 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U81 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U82 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U30 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U29 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U30 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U298 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0048 * d[1])))) + (16'(16'h0018 * d[2])))) + (16'(16'h0008 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U297 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U298 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0002;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U275 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U274 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U275 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U252 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U251 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U252 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U229 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001c * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U228 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [2:0];
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U229 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_next_value_out = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U177 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0984 * d[1])))) + (16'(16'h032c * d[2])))) + (16'(16'h001d * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U176 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire d_4_at_max_out;
wire [15:0] d_4_next_value_out;
wire [15:0] d_4_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [4:0];
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U177 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_next_value_out = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_next_value_out = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_next_value_out),
    .clk(clk),
    .out(d_4_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U134 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0310 * d[1])))) + (16'(16'h001c * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h3e91);
endmodule

module affine_controller__U133 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [3:0];
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U134 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_next_value_out = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_next_value_out = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_next_value_out = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h00f0 * d[1])))) + (16'(16'h0008 * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h0001);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire cmp_time_out;
wire [15:0] cycle_time_out;
wire [15:0] d_0_next_value_out;
wire [15:0] d_0_reg_out;
wire d_1_at_max_out;
wire [15:0] d_1_next_value_out;
wire [15:0] d_1_reg_out;
wire d_2_at_max_out;
wire [15:0] d_2_next_value_out;
wire [15:0] d_2_reg_out;
wire d_3_at_max_out;
wire [15:0] d_3_next_value_out;
wire [15:0] d_3_reg_out;
wire [15:0] inc_time_out;
wire [15:0] affine_func_d [3:0];
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(inc_time_out),
    .clk(clk),
    .out(cycle_time_out)
);
assign d_0_next_value_out = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_next_value_out),
    .clk(clk),
    .out(d_0_reg_out),
    .en(cmp_time_out)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_next_value_out = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_next_value_out),
    .clk(clk),
    .out(d_1_reg_out),
    .en(cmp_time_out)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_next_value_out = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_next_value_out),
    .clk(clk),
    .out(d_2_reg_out),
    .en(cmp_time_out)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_next_value_out = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_next_value_out),
    .clk(clk),
    .out(d_3_reg_out),
    .en(cmp_time_out)
);
assign inc_time_out = 16'(cycle_time_out + 16'h0001);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] arr__U116_out [4:0];
wire [15:0] arr__U126_out [4:0];
wire [15:0] arr__U161_out [3:0];
wire [15:0] arr__U170_out [3:0];
wire [15:0] arr__U211_out [4:0];
wire [15:0] arr__U221_out [4:0];
wire [15:0] arr__U64_out [4:0];
wire [15:0] arr__U74_out [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U114_out;
wire delay_reg__U124_out;
wire delay_reg__U159_out;
wire delay_reg__U168_out;
wire delay_reg__U209_out;
wire delay_reg__U219_out;
wire delay_reg__U62_out;
wire delay_reg__U72_out;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
wire [15:0] arr__U116_in [4:0];
assign arr__U116_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U116_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U116_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U116_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U116_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U117 arr__U116 (
    .clk(clk),
    .in(arr__U116_in),
    .out(arr__U116_out)
);
wire [15:0] arr__U126_in [4:0];
assign arr__U126_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U126_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U126_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U126_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U126_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U127 arr__U126 (
    .clk(clk),
    .in(arr__U126_in),
    .out(arr__U126_out)
);
wire [15:0] arr__U161_in [3:0];
assign arr__U161_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U161_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U161_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U161_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U162 arr__U161 (
    .clk(clk),
    .in(arr__U161_in),
    .out(arr__U161_out)
);
wire [15:0] arr__U170_in [3:0];
assign arr__U170_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U170_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U170_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U170_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U171 arr__U170 (
    .clk(clk),
    .in(arr__U170_in),
    .out(arr__U170_out)
);
wire [15:0] arr__U211_in [4:0];
assign arr__U211_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U211_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U211_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U211_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U211_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U212 arr__U211 (
    .clk(clk),
    .in(arr__U211_in),
    .out(arr__U211_out)
);
wire [15:0] arr__U221_in [4:0];
assign arr__U221_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U221_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U221_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U221_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U221_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U222 arr__U221 (
    .clk(clk),
    .in(arr__U221_in),
    .out(arr__U221_out)
);
wire [15:0] arr__U64_in [4:0];
assign arr__U64_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U64_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U64_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U64_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U64_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U65 arr__U64 (
    .clk(clk),
    .in(arr__U64_in),
    .out(arr__U64_out)
);
wire [15:0] arr__U74_in [4:0];
assign arr__U74_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U74_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U74_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U74_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U74_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U75 arr__U74 (
    .clk(clk),
    .in(arr__U74_in),
    .out(arr__U74_out)
);
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_1_write_wen(op_hcompute_conv_stencil_1_write_start_out),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(op_hcompute_conv_stencil_2_write_start_out),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(op_hcompute_conv_stencil_3_read_start_out),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(op_hcompute_conv_stencil_3_write_start_out),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(op_hcompute_conv_stencil_4_read_start_out),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(op_hcompute_conv_stencil_4_write_start_out),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(op_hcompute_conv_stencil_5_read_start_out),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(op_hcompute_conv_stencil_5_write_start_out),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(op_hcompute_conv_stencil_write_start_out),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(op_hcompute_hw_output_stencil_read_start_out),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U114 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(delay_reg__U114_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U124 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(delay_reg__U124_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U159 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(delay_reg__U159_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U168 (
    .clk(clk),
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(delay_reg__U168_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U209 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(delay_reg__U209_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U219 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(delay_reg__U219_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U62 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(delay_reg__U62_out)
);
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U72 (
    .clk(clk),
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(delay_reg__U72_out)
);
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_3_read_ren(op_hcompute_conv_stencil_3_read_start_out),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(op_hcompute_conv_stencil_4_read_start_out),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(op_hcompute_conv_stencil_5_read_start_out),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(op_hcompute_hw_input_global_wrapper_stencil_write_start_out),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(clk),
    .flush(flush),
    .rst_n(rst_n),
    .op_hcompute_conv_stencil_3_read_ren(op_hcompute_conv_stencil_3_read_start_out),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(op_hcompute_conv_stencil_4_read_start_out),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(op_hcompute_conv_stencil_5_read_start_out),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
op_hcompute_conv_stencil_1_exe_start_pt__U270 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U271 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
affine_controller__U251 op_hcompute_conv_stencil_1_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
op_hcompute_conv_stencil_1_read_start_pt__U268 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U269 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
op_hcompute_conv_stencil_1_write_start_pt__U272 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_port_controller_valid),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U273 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
op_hcompute_conv_stencil_2_exe_start_pt__U247 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U248 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
affine_controller__U228 op_hcompute_conv_stencil_2_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
op_hcompute_conv_stencil_2_read_start_pt__U245 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U246 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
op_hcompute_conv_stencil_2_write_start_pt__U249 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_port_controller_valid),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U250 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
op_hcompute_conv_stencil_3_exe_start_pt__U113 op_hcompute_conv_stencil_3_exe_start (
    .in(delay_reg__U114_out),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U116_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U116_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U116_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U116_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U116_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U115 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
affine_controller__U81 op_hcompute_conv_stencil_3_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
op_hcompute_conv_stencil_3_read_start_pt__U111 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_port_controller_valid),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U112 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
op_hcompute_conv_stencil_3_write_start_pt__U123 op_hcompute_conv_stencil_3_write_start (
    .in(delay_reg__U124_out),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U126_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U126_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U126_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U126_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U126_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U125 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
op_hcompute_conv_stencil_4_exe_start_pt__U61 op_hcompute_conv_stencil_4_exe_start (
    .in(delay_reg__U62_out),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U64_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U64_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U64_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U64_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U64_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U63 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
affine_controller__U29 op_hcompute_conv_stencil_4_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
op_hcompute_conv_stencil_4_read_start_pt__U59 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_port_controller_valid),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U60 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
op_hcompute_conv_stencil_4_write_start_pt__U71 op_hcompute_conv_stencil_4_write_start (
    .in(delay_reg__U72_out),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U74_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U74_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U74_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U74_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U74_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U73 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
op_hcompute_conv_stencil_5_exe_start_pt__U208 op_hcompute_conv_stencil_5_exe_start (
    .in(delay_reg__U209_out),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U211_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U211_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U211_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U211_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U211_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U210 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
affine_controller__U176 op_hcompute_conv_stencil_5_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
op_hcompute_conv_stencil_5_read_start_pt__U206 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_port_controller_valid),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U207 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
op_hcompute_conv_stencil_5_write_start_pt__U218 op_hcompute_conv_stencil_5_write_start (
    .in(delay_reg__U219_out),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U221_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U221_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U221_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U221_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U221_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U220 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
op_hcompute_conv_stencil_exe_start_pt__U293 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U294 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
affine_controller__U274 op_hcompute_conv_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
op_hcompute_conv_stencil_read_start_pt__U291 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_read_start_out)
);
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U292 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
op_hcompute_conv_stencil_write_start_pt__U295 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_port_controller_valid),
    .out(op_hcompute_conv_stencil_write_start_out)
);
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U296 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U25 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U26 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
affine_controller__U0 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U23 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U24 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U27 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U28 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U329 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U330 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
affine_controller__U297 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U327 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U328 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U331 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U332 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
op_hcompute_hw_output_stencil_exe_start_pt__U158 op_hcompute_hw_output_stencil_exe_start (
    .in(delay_reg__U159_out),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U161_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U161_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U161_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U161_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U160 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
affine_controller__U133 op_hcompute_hw_output_stencil_port_controller (
    .clk(clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
op_hcompute_hw_output_stencil_read_start_pt__U156 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_port_controller_valid),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U157 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
op_hcompute_hw_output_stencil_write_start_pt__U167 op_hcompute_hw_output_stencil_write_start (
    .in(delay_reg__U168_out),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U170_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U170_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U170_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U170_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U169 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

