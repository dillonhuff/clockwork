// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U739 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U742 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U721 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U722 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U723 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U726 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U696 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U697 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U692 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U693 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U694 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U695 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U27 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U28 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U23 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U24 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U25 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U26 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U261 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U262 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U257 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U258 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U259 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U260 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U313 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U331 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U293 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U294 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U295 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U298 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U102 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U120 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U82 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U83 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U84 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U87 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U524 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U542 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U504 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U505 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U506 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U509 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U472 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U473 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U468 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U469 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U470 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U471 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U50 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U51 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U46 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U47 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U48 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U49 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U96 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U97_in;
wire _U97_clk;
wire [15:0] _U97_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U100_in = in[3];
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = in[4];
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U97_in = in[0];
assign _U97_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(_U97_in),
    .clk(_U97_clk),
    .out(_U97_out)
);
assign _U98_in = in[1];
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = in[2];
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
assign out[4] = _U101_out;
assign out[3] = _U100_out;
assign out[2] = _U99_out;
assign out[1] = _U98_out;
assign out[0] = _U97_out;
endmodule

module array_delay_U89 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
wire [15:0] _U93_in;
wire _U93_clk;
wire [15:0] _U93_out;
wire [15:0] _U94_in;
wire _U94_clk;
wire [15:0] _U94_out;
assign _U90_in = in[0];
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = in[1];
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = in[2];
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign _U93_in = in[3];
assign _U93_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U93_in),
    .clk(_U93_clk),
    .out(_U93_out)
);
assign _U94_in = in[4];
assign _U94_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U94_in),
    .clk(_U94_clk),
    .out(_U94_out)
);
assign out[4] = _U94_out;
assign out[3] = _U93_out;
assign out[2] = _U92_out;
assign out[1] = _U91_out;
assign out[0] = _U90_out;
endmodule

module array_delay_U750 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U751_in;
wire _U751_clk;
wire [15:0] _U751_out;
wire [15:0] _U752_in;
wire _U752_clk;
wire [15:0] _U752_out;
wire [15:0] _U753_in;
wire _U753_clk;
wire [15:0] _U753_out;
wire [15:0] _U754_in;
wire _U754_clk;
wire [15:0] _U754_out;
assign _U751_in = in[0];
assign _U751_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U751 (
    .in(_U751_in),
    .clk(_U751_clk),
    .out(_U751_out)
);
assign _U752_in = in[1];
assign _U752_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U752 (
    .in(_U752_in),
    .clk(_U752_clk),
    .out(_U752_out)
);
assign _U753_in = in[2];
assign _U753_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U753 (
    .in(_U753_in),
    .clk(_U753_clk),
    .out(_U753_out)
);
assign _U754_in = in[3];
assign _U754_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U754 (
    .in(_U754_in),
    .clk(_U754_clk),
    .out(_U754_out)
);
assign out[3] = _U754_out;
assign out[2] = _U753_out;
assign out[1] = _U752_out;
assign out[0] = _U751_out;
endmodule

module array_delay_U744 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U745_in;
wire _U745_clk;
wire [15:0] _U745_out;
wire [15:0] _U746_in;
wire _U746_clk;
wire [15:0] _U746_out;
wire [15:0] _U747_in;
wire _U747_clk;
wire [15:0] _U747_out;
wire [15:0] _U748_in;
wire _U748_clk;
wire [15:0] _U748_out;
assign _U745_in = in[0];
assign _U745_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U745 (
    .in(_U745_in),
    .clk(_U745_clk),
    .out(_U745_out)
);
assign _U746_in = in[1];
assign _U746_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U746 (
    .in(_U746_in),
    .clk(_U746_clk),
    .out(_U746_out)
);
assign _U747_in = in[2];
assign _U747_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U747 (
    .in(_U747_in),
    .clk(_U747_clk),
    .out(_U747_out)
);
assign _U748_in = in[3];
assign _U748_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U748 (
    .in(_U748_in),
    .clk(_U748_clk),
    .out(_U748_out)
);
assign out[3] = _U748_out;
assign out[2] = _U747_out;
assign out[1] = _U746_out;
assign out[0] = _U745_out;
endmodule

module array_delay_U734 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U735_in;
wire _U735_clk;
wire [15:0] _U735_out;
wire [15:0] _U736_in;
wire _U736_clk;
wire [15:0] _U736_out;
wire [15:0] _U737_in;
wire _U737_clk;
wire [15:0] _U737_out;
wire [15:0] _U738_in;
wire _U738_clk;
wire [15:0] _U738_out;
assign _U735_in = in[0];
assign _U735_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U735 (
    .in(_U735_in),
    .clk(_U735_clk),
    .out(_U735_out)
);
assign _U736_in = in[1];
assign _U736_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U736 (
    .in(_U736_in),
    .clk(_U736_clk),
    .out(_U736_out)
);
assign _U737_in = in[2];
assign _U737_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U737 (
    .in(_U737_in),
    .clk(_U737_clk),
    .out(_U737_out)
);
assign _U738_in = in[3];
assign _U738_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U738 (
    .in(_U738_in),
    .clk(_U738_clk),
    .out(_U738_out)
);
assign out[3] = _U738_out;
assign out[2] = _U737_out;
assign out[1] = _U736_out;
assign out[0] = _U735_out;
endmodule

module array_delay_U728 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U729_in;
wire _U729_clk;
wire [15:0] _U729_out;
wire [15:0] _U730_in;
wire _U730_clk;
wire [15:0] _U730_out;
wire [15:0] _U731_in;
wire _U731_clk;
wire [15:0] _U731_out;
wire [15:0] _U732_in;
wire _U732_clk;
wire [15:0] _U732_out;
assign _U729_in = in[0];
assign _U729_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U729 (
    .in(_U729_in),
    .clk(_U729_clk),
    .out(_U729_out)
);
assign _U730_in = in[1];
assign _U730_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U730 (
    .in(_U730_in),
    .clk(_U730_clk),
    .out(_U730_out)
);
assign _U731_in = in[2];
assign _U731_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U731 (
    .in(_U731_in),
    .clk(_U731_clk),
    .out(_U731_out)
);
assign _U732_in = in[3];
assign _U732_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U732 (
    .in(_U732_in),
    .clk(_U732_clk),
    .out(_U732_out)
);
assign out[3] = _U732_out;
assign out[2] = _U731_out;
assign out[1] = _U730_out;
assign out[0] = _U729_out;
endmodule

module array_delay_U656 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U657_in;
wire _U657_clk;
wire [15:0] _U657_out;
wire [15:0] _U658_in;
wire _U658_clk;
wire [15:0] _U658_out;
wire [15:0] _U659_in;
wire _U659_clk;
wire [15:0] _U659_out;
wire [15:0] _U660_in;
wire _U660_clk;
wire [15:0] _U660_out;
wire [15:0] _U661_in;
wire _U661_clk;
wire [15:0] _U661_out;
assign _U657_in = in[0];
assign _U657_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U657 (
    .in(_U657_in),
    .clk(_U657_clk),
    .out(_U657_out)
);
assign _U658_in = in[1];
assign _U658_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U658 (
    .in(_U658_in),
    .clk(_U658_clk),
    .out(_U658_out)
);
assign _U659_in = in[2];
assign _U659_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U659 (
    .in(_U659_in),
    .clk(_U659_clk),
    .out(_U659_out)
);
assign _U660_in = in[3];
assign _U660_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U660 (
    .in(_U660_in),
    .clk(_U660_clk),
    .out(_U660_out)
);
assign _U661_in = in[4];
assign _U661_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U661 (
    .in(_U661_in),
    .clk(_U661_clk),
    .out(_U661_out)
);
assign out[4] = _U661_out;
assign out[3] = _U660_out;
assign out[2] = _U659_out;
assign out[1] = _U658_out;
assign out[0] = _U657_out;
endmodule

module array_delay_U649 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U650_in;
wire _U650_clk;
wire [15:0] _U650_out;
wire [15:0] _U651_in;
wire _U651_clk;
wire [15:0] _U651_out;
wire [15:0] _U652_in;
wire _U652_clk;
wire [15:0] _U652_out;
wire [15:0] _U653_in;
wire _U653_clk;
wire [15:0] _U653_out;
wire [15:0] _U654_in;
wire _U654_clk;
wire [15:0] _U654_out;
assign _U650_in = in[0];
assign _U650_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U650 (
    .in(_U650_in),
    .clk(_U650_clk),
    .out(_U650_out)
);
assign _U651_in = in[1];
assign _U651_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U651 (
    .in(_U651_in),
    .clk(_U651_clk),
    .out(_U651_out)
);
assign _U652_in = in[2];
assign _U652_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U652 (
    .in(_U652_in),
    .clk(_U652_clk),
    .out(_U652_out)
);
assign _U653_in = in[3];
assign _U653_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U653 (
    .in(_U653_in),
    .clk(_U653_clk),
    .out(_U653_out)
);
assign _U654_in = in[4];
assign _U654_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U654 (
    .in(_U654_in),
    .clk(_U654_clk),
    .out(_U654_out)
);
assign out[4] = _U654_out;
assign out[3] = _U653_out;
assign out[2] = _U652_out;
assign out[1] = _U651_out;
assign out[0] = _U650_out;
endmodule

module array_delay_U642 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U643_in;
wire _U643_clk;
wire [15:0] _U643_out;
wire [15:0] _U644_in;
wire _U644_clk;
wire [15:0] _U644_out;
wire [15:0] _U645_in;
wire _U645_clk;
wire [15:0] _U645_out;
wire [15:0] _U646_in;
wire _U646_clk;
wire [15:0] _U646_out;
wire [15:0] _U647_in;
wire _U647_clk;
wire [15:0] _U647_out;
assign _U643_in = in[0];
assign _U643_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U643 (
    .in(_U643_in),
    .clk(_U643_clk),
    .out(_U643_out)
);
assign _U644_in = in[1];
assign _U644_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U644 (
    .in(_U644_in),
    .clk(_U644_clk),
    .out(_U644_out)
);
assign _U645_in = in[2];
assign _U645_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U645 (
    .in(_U645_in),
    .clk(_U645_clk),
    .out(_U645_out)
);
assign _U646_in = in[3];
assign _U646_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U646 (
    .in(_U646_in),
    .clk(_U646_clk),
    .out(_U646_out)
);
assign _U647_in = in[4];
assign _U647_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U647 (
    .in(_U647_in),
    .clk(_U647_clk),
    .out(_U647_out)
);
assign out[4] = _U647_out;
assign out[3] = _U646_out;
assign out[2] = _U645_out;
assign out[1] = _U644_out;
assign out[0] = _U643_out;
endmodule

module array_delay_U635 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U636_in;
wire _U636_clk;
wire [15:0] _U636_out;
wire [15:0] _U637_in;
wire _U637_clk;
wire [15:0] _U637_out;
wire [15:0] _U638_in;
wire _U638_clk;
wire [15:0] _U638_out;
wire [15:0] _U639_in;
wire _U639_clk;
wire [15:0] _U639_out;
wire [15:0] _U640_in;
wire _U640_clk;
wire [15:0] _U640_out;
assign _U636_in = in[0];
assign _U636_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U636 (
    .in(_U636_in),
    .clk(_U636_clk),
    .out(_U636_out)
);
assign _U637_in = in[1];
assign _U637_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U637 (
    .in(_U637_in),
    .clk(_U637_clk),
    .out(_U637_out)
);
assign _U638_in = in[2];
assign _U638_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U638 (
    .in(_U638_in),
    .clk(_U638_clk),
    .out(_U638_out)
);
assign _U639_in = in[3];
assign _U639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(_U639_in),
    .clk(_U639_clk),
    .out(_U639_out)
);
assign _U640_in = in[4];
assign _U640_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U640 (
    .in(_U640_in),
    .clk(_U640_clk),
    .out(_U640_out)
);
assign out[4] = _U640_out;
assign out[3] = _U639_out;
assign out[2] = _U638_out;
assign out[1] = _U637_out;
assign out[0] = _U636_out;
endmodule

module array_delay_U628 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U629_in;
wire _U629_clk;
wire [15:0] _U629_out;
wire [15:0] _U630_in;
wire _U630_clk;
wire [15:0] _U630_out;
wire [15:0] _U631_in;
wire _U631_clk;
wire [15:0] _U631_out;
wire [15:0] _U632_in;
wire _U632_clk;
wire [15:0] _U632_out;
wire [15:0] _U633_in;
wire _U633_clk;
wire [15:0] _U633_out;
assign _U629_in = in[0];
assign _U629_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U629 (
    .in(_U629_in),
    .clk(_U629_clk),
    .out(_U629_out)
);
assign _U630_in = in[1];
assign _U630_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U630 (
    .in(_U630_in),
    .clk(_U630_clk),
    .out(_U630_out)
);
assign _U631_in = in[2];
assign _U631_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U631 (
    .in(_U631_in),
    .clk(_U631_clk),
    .out(_U631_out)
);
assign _U632_in = in[3];
assign _U632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(_U632_in),
    .clk(_U632_clk),
    .out(_U632_out)
);
assign _U633_in = in[4];
assign _U633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(_U633_in),
    .clk(_U633_clk),
    .out(_U633_out)
);
assign out[4] = _U633_out;
assign out[3] = _U632_out;
assign out[2] = _U631_out;
assign out[1] = _U630_out;
assign out[0] = _U629_out;
endmodule

module array_delay_U621 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U622_in;
wire _U622_clk;
wire [15:0] _U622_out;
wire [15:0] _U623_in;
wire _U623_clk;
wire [15:0] _U623_out;
wire [15:0] _U624_in;
wire _U624_clk;
wire [15:0] _U624_out;
wire [15:0] _U625_in;
wire _U625_clk;
wire [15:0] _U625_out;
wire [15:0] _U626_in;
wire _U626_clk;
wire [15:0] _U626_out;
assign _U622_in = in[0];
assign _U622_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U622 (
    .in(_U622_in),
    .clk(_U622_clk),
    .out(_U622_out)
);
assign _U623_in = in[1];
assign _U623_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U623 (
    .in(_U623_in),
    .clk(_U623_clk),
    .out(_U623_out)
);
assign _U624_in = in[2];
assign _U624_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U624 (
    .in(_U624_in),
    .clk(_U624_clk),
    .out(_U624_out)
);
assign _U625_in = in[3];
assign _U625_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U625 (
    .in(_U625_in),
    .clk(_U625_clk),
    .out(_U625_out)
);
assign _U626_in = in[4];
assign _U626_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U626 (
    .in(_U626_in),
    .clk(_U626_clk),
    .out(_U626_out)
);
assign out[4] = _U626_out;
assign out[3] = _U625_out;
assign out[2] = _U624_out;
assign out[1] = _U623_out;
assign out[0] = _U622_out;
endmodule

module array_delay_U614 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U615_in;
wire _U615_clk;
wire [15:0] _U615_out;
wire [15:0] _U616_in;
wire _U616_clk;
wire [15:0] _U616_out;
wire [15:0] _U617_in;
wire _U617_clk;
wire [15:0] _U617_out;
wire [15:0] _U618_in;
wire _U618_clk;
wire [15:0] _U618_out;
wire [15:0] _U619_in;
wire _U619_clk;
wire [15:0] _U619_out;
assign _U615_in = in[0];
assign _U615_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U615 (
    .in(_U615_in),
    .clk(_U615_clk),
    .out(_U615_out)
);
assign _U616_in = in[1];
assign _U616_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U616 (
    .in(_U616_in),
    .clk(_U616_clk),
    .out(_U616_out)
);
assign _U617_in = in[2];
assign _U617_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U617 (
    .in(_U617_in),
    .clk(_U617_clk),
    .out(_U617_out)
);
assign _U618_in = in[3];
assign _U618_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U618 (
    .in(_U618_in),
    .clk(_U618_clk),
    .out(_U618_out)
);
assign _U619_in = in[4];
assign _U619_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U619 (
    .in(_U619_in),
    .clk(_U619_clk),
    .out(_U619_out)
);
assign out[4] = _U619_out;
assign out[3] = _U618_out;
assign out[2] = _U617_out;
assign out[1] = _U616_out;
assign out[0] = _U615_out;
endmodule

module array_delay_U607 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U608_in;
wire _U608_clk;
wire [15:0] _U608_out;
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
wire [15:0] _U611_in;
wire _U611_clk;
wire [15:0] _U611_out;
wire [15:0] _U612_in;
wire _U612_clk;
wire [15:0] _U612_out;
assign _U608_in = in[0];
assign _U608_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U608 (
    .in(_U608_in),
    .clk(_U608_clk),
    .out(_U608_out)
);
assign _U609_in = in[1];
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = in[2];
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
assign _U611_in = in[3];
assign _U611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U611 (
    .in(_U611_in),
    .clk(_U611_clk),
    .out(_U611_out)
);
assign _U612_in = in[4];
assign _U612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U612 (
    .in(_U612_in),
    .clk(_U612_clk),
    .out(_U612_out)
);
assign out[4] = _U612_out;
assign out[3] = _U611_out;
assign out[2] = _U610_out;
assign out[1] = _U609_out;
assign out[0] = _U608_out;
endmodule

module array_delay_U600 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U601_in;
wire _U601_clk;
wire [15:0] _U601_out;
wire [15:0] _U602_in;
wire _U602_clk;
wire [15:0] _U602_out;
wire [15:0] _U603_in;
wire _U603_clk;
wire [15:0] _U603_out;
wire [15:0] _U604_in;
wire _U604_clk;
wire [15:0] _U604_out;
wire [15:0] _U605_in;
wire _U605_clk;
wire [15:0] _U605_out;
assign _U601_in = in[0];
assign _U601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U601_in),
    .clk(_U601_clk),
    .out(_U601_out)
);
assign _U602_in = in[1];
assign _U602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U602_in),
    .clk(_U602_clk),
    .out(_U602_out)
);
assign _U603_in = in[2];
assign _U603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U603 (
    .in(_U603_in),
    .clk(_U603_clk),
    .out(_U603_out)
);
assign _U604_in = in[3];
assign _U604_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U604 (
    .in(_U604_in),
    .clk(_U604_clk),
    .out(_U604_out)
);
assign _U605_in = in[4];
assign _U605_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U605 (
    .in(_U605_in),
    .clk(_U605_clk),
    .out(_U605_out)
);
assign out[4] = _U605_out;
assign out[3] = _U604_out;
assign out[2] = _U603_out;
assign out[1] = _U602_out;
assign out[0] = _U601_out;
endmodule

module array_delay_U593 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U594_in;
wire _U594_clk;
wire [15:0] _U594_out;
wire [15:0] _U595_in;
wire _U595_clk;
wire [15:0] _U595_out;
wire [15:0] _U596_in;
wire _U596_clk;
wire [15:0] _U596_out;
wire [15:0] _U597_in;
wire _U597_clk;
wire [15:0] _U597_out;
wire [15:0] _U598_in;
wire _U598_clk;
wire [15:0] _U598_out;
assign _U594_in = in[0];
assign _U594_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U594 (
    .in(_U594_in),
    .clk(_U594_clk),
    .out(_U594_out)
);
assign _U595_in = in[1];
assign _U595_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U595 (
    .in(_U595_in),
    .clk(_U595_clk),
    .out(_U595_out)
);
assign _U596_in = in[2];
assign _U596_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U596 (
    .in(_U596_in),
    .clk(_U596_clk),
    .out(_U596_out)
);
assign _U597_in = in[3];
assign _U597_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U597 (
    .in(_U597_in),
    .clk(_U597_clk),
    .out(_U597_out)
);
assign _U598_in = in[4];
assign _U598_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U598 (
    .in(_U598_in),
    .clk(_U598_clk),
    .out(_U598_out)
);
assign out[4] = _U598_out;
assign out[3] = _U597_out;
assign out[2] = _U596_out;
assign out[1] = _U595_out;
assign out[0] = _U594_out;
endmodule

module array_delay_U586 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U587_in;
wire _U587_clk;
wire [15:0] _U587_out;
wire [15:0] _U588_in;
wire _U588_clk;
wire [15:0] _U588_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
assign _U587_in = in[0];
assign _U587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U587_in),
    .clk(_U587_clk),
    .out(_U587_out)
);
assign _U588_in = in[1];
assign _U588_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(_U588_in),
    .clk(_U588_clk),
    .out(_U588_out)
);
assign _U589_in = in[2];
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = in[3];
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = in[4];
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign out[4] = _U591_out;
assign out[3] = _U590_out;
assign out[2] = _U589_out;
assign out[1] = _U588_out;
assign out[0] = _U587_out;
endmodule

module array_delay_U579 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U580_in;
wire _U580_clk;
wire [15:0] _U580_out;
wire [15:0] _U581_in;
wire _U581_clk;
wire [15:0] _U581_out;
wire [15:0] _U582_in;
wire _U582_clk;
wire [15:0] _U582_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
assign _U580_in = in[0];
assign _U580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U580_in),
    .clk(_U580_clk),
    .out(_U580_out)
);
assign _U581_in = in[1];
assign _U581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U581_in),
    .clk(_U581_clk),
    .out(_U581_out)
);
assign _U582_in = in[2];
assign _U582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U582_in),
    .clk(_U582_clk),
    .out(_U582_out)
);
assign _U583_in = in[3];
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = in[4];
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign out[4] = _U584_out;
assign out[3] = _U583_out;
assign out[2] = _U582_out;
assign out[1] = _U581_out;
assign out[0] = _U580_out;
endmodule

module array_delay_U572 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U573_in;
wire _U573_clk;
wire [15:0] _U573_out;
wire [15:0] _U574_in;
wire _U574_clk;
wire [15:0] _U574_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire _U576_clk;
wire [15:0] _U576_out;
wire [15:0] _U577_in;
wire _U577_clk;
wire [15:0] _U577_out;
assign _U573_in = in[0];
assign _U573_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U573 (
    .in(_U573_in),
    .clk(_U573_clk),
    .out(_U573_out)
);
assign _U574_in = in[1];
assign _U574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(_U574_in),
    .clk(_U574_clk),
    .out(_U574_out)
);
assign _U575_in = in[2];
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = in[3];
assign _U576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U576_in),
    .clk(_U576_clk),
    .out(_U576_out)
);
assign _U577_in = in[4];
assign _U577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U577 (
    .in(_U577_in),
    .clk(_U577_clk),
    .out(_U577_out)
);
assign out[4] = _U577_out;
assign out[3] = _U576_out;
assign out[2] = _U575_out;
assign out[1] = _U574_out;
assign out[0] = _U573_out;
endmodule

module array_delay_U565 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U566_in;
wire _U566_clk;
wire [15:0] _U566_out;
wire [15:0] _U567_in;
wire _U567_clk;
wire [15:0] _U567_out;
wire [15:0] _U568_in;
wire _U568_clk;
wire [15:0] _U568_out;
wire [15:0] _U569_in;
wire _U569_clk;
wire [15:0] _U569_out;
wire [15:0] _U570_in;
wire _U570_clk;
wire [15:0] _U570_out;
assign _U566_in = in[0];
assign _U566_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(_U566_in),
    .clk(_U566_clk),
    .out(_U566_out)
);
assign _U567_in = in[1];
assign _U567_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U567 (
    .in(_U567_in),
    .clk(_U567_clk),
    .out(_U567_out)
);
assign _U568_in = in[2];
assign _U568_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U568 (
    .in(_U568_in),
    .clk(_U568_clk),
    .out(_U568_out)
);
assign _U569_in = in[3];
assign _U569_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(_U569_in),
    .clk(_U569_clk),
    .out(_U569_out)
);
assign _U570_in = in[4];
assign _U570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U570_in),
    .clk(_U570_clk),
    .out(_U570_out)
);
assign out[4] = _U570_out;
assign out[3] = _U569_out;
assign out[2] = _U568_out;
assign out[1] = _U567_out;
assign out[0] = _U566_out;
endmodule

module array_delay_U558 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U559_in;
wire _U559_clk;
wire [15:0] _U559_out;
wire [15:0] _U560_in;
wire _U560_clk;
wire [15:0] _U560_out;
wire [15:0] _U561_in;
wire _U561_clk;
wire [15:0] _U561_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
assign _U559_in = in[0];
assign _U559_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U559 (
    .in(_U559_in),
    .clk(_U559_clk),
    .out(_U559_out)
);
assign _U560_in = in[1];
assign _U560_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U560 (
    .in(_U560_in),
    .clk(_U560_clk),
    .out(_U560_out)
);
assign _U561_in = in[2];
assign _U561_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(_U561_in),
    .clk(_U561_clk),
    .out(_U561_out)
);
assign _U562_in = in[3];
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = in[4];
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign out[4] = _U563_out;
assign out[3] = _U562_out;
assign out[2] = _U561_out;
assign out[1] = _U560_out;
assign out[0] = _U559_out;
endmodule

module array_delay_U551 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire _U553_clk;
wire [15:0] _U553_out;
wire [15:0] _U554_in;
wire _U554_clk;
wire [15:0] _U554_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
assign _U552_in = in[0];
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = in[1];
assign _U553_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U553 (
    .in(_U553_in),
    .clk(_U553_clk),
    .out(_U553_out)
);
assign _U554_in = in[2];
assign _U554_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U554 (
    .in(_U554_in),
    .clk(_U554_clk),
    .out(_U554_out)
);
assign _U555_in = in[3];
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = in[4];
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign out[4] = _U556_out;
assign out[3] = _U555_out;
assign out[2] = _U554_out;
assign out[1] = _U553_out;
assign out[0] = _U552_out;
endmodule

module array_delay_U544 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
wire [15:0] _U547_in;
wire _U547_clk;
wire [15:0] _U547_out;
wire [15:0] _U548_in;
wire _U548_clk;
wire [15:0] _U548_out;
wire [15:0] _U549_in;
wire _U549_clk;
wire [15:0] _U549_out;
assign _U545_in = in[0];
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = in[1];
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign _U547_in = in[2];
assign _U547_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(_U547_in),
    .clk(_U547_clk),
    .out(_U547_out)
);
assign _U548_in = in[3];
assign _U548_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(_U548_in),
    .clk(_U548_clk),
    .out(_U548_out)
);
assign _U549_in = in[4];
assign _U549_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U549 (
    .in(_U549_in),
    .clk(_U549_clk),
    .out(_U549_out)
);
assign out[4] = _U549_out;
assign out[3] = _U548_out;
assign out[2] = _U547_out;
assign out[1] = _U546_out;
assign out[0] = _U545_out;
endmodule

module array_delay_U518 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire _U520_clk;
wire [15:0] _U520_out;
wire [15:0] _U521_in;
wire _U521_clk;
wire [15:0] _U521_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
assign _U519_in = in[0];
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = in[1];
assign _U520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U520_in),
    .clk(_U520_clk),
    .out(_U520_out)
);
assign _U521_in = in[2];
assign _U521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U521_in),
    .clk(_U521_clk),
    .out(_U521_out)
);
assign _U522_in = in[3];
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = in[4];
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign out[4] = _U523_out;
assign out[3] = _U522_out;
assign out[2] = _U521_out;
assign out[1] = _U520_out;
assign out[0] = _U519_out;
endmodule

module array_delay_U511 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire _U513_clk;
wire [15:0] _U513_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
assign _U512_in = in[0];
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = in[1];
assign _U513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U513_in),
    .clk(_U513_clk),
    .out(_U513_out)
);
assign _U514_in = in[2];
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = in[3];
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = in[4];
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign out[4] = _U516_out;
assign out[3] = _U515_out;
assign out[2] = _U514_out;
assign out[1] = _U513_out;
assign out[0] = _U512_out;
endmodule

module array_delay_U445 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
wire [15:0] _U447_in;
wire _U447_clk;
wire [15:0] _U447_out;
wire [15:0] _U448_in;
wire _U448_clk;
wire [15:0] _U448_out;
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
assign _U446_in = in[0];
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign _U447_in = in[1];
assign _U447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U447 (
    .in(_U447_in),
    .clk(_U447_clk),
    .out(_U447_out)
);
assign _U448_in = in[2];
assign _U448_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U448 (
    .in(_U448_in),
    .clk(_U448_clk),
    .out(_U448_out)
);
assign _U449_in = in[3];
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = in[4];
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign out[4] = _U450_out;
assign out[3] = _U449_out;
assign out[2] = _U448_out;
assign out[1] = _U447_out;
assign out[0] = _U446_out;
endmodule

module array_delay_U438 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
assign _U439_in = in[0];
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign _U440_in = in[1];
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = in[2];
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign _U442_in = in[3];
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = in[4];
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign out[4] = _U443_out;
assign out[3] = _U442_out;
assign out[2] = _U441_out;
assign out[1] = _U440_out;
assign out[0] = _U439_out;
endmodule

module array_delay_U431 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U432_in;
wire _U432_clk;
wire [15:0] _U432_out;
wire [15:0] _U433_in;
wire _U433_clk;
wire [15:0] _U433_out;
wire [15:0] _U434_in;
wire _U434_clk;
wire [15:0] _U434_out;
wire [15:0] _U435_in;
wire _U435_clk;
wire [15:0] _U435_out;
wire [15:0] _U436_in;
wire _U436_clk;
wire [15:0] _U436_out;
assign _U432_in = in[0];
assign _U432_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U432 (
    .in(_U432_in),
    .clk(_U432_clk),
    .out(_U432_out)
);
assign _U433_in = in[1];
assign _U433_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U433 (
    .in(_U433_in),
    .clk(_U433_clk),
    .out(_U433_out)
);
assign _U434_in = in[2];
assign _U434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U434_in),
    .clk(_U434_clk),
    .out(_U434_out)
);
assign _U435_in = in[3];
assign _U435_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U435 (
    .in(_U435_in),
    .clk(_U435_clk),
    .out(_U435_out)
);
assign _U436_in = in[4];
assign _U436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U436 (
    .in(_U436_in),
    .clk(_U436_clk),
    .out(_U436_out)
);
assign out[4] = _U436_out;
assign out[3] = _U435_out;
assign out[2] = _U434_out;
assign out[1] = _U433_out;
assign out[0] = _U432_out;
endmodule

module array_delay_U424 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U425_in;
wire _U425_clk;
wire [15:0] _U425_out;
wire [15:0] _U426_in;
wire _U426_clk;
wire [15:0] _U426_out;
wire [15:0] _U427_in;
wire _U427_clk;
wire [15:0] _U427_out;
wire [15:0] _U428_in;
wire _U428_clk;
wire [15:0] _U428_out;
wire [15:0] _U429_in;
wire _U429_clk;
wire [15:0] _U429_out;
assign _U425_in = in[0];
assign _U425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U425 (
    .in(_U425_in),
    .clk(_U425_clk),
    .out(_U425_out)
);
assign _U426_in = in[1];
assign _U426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U426 (
    .in(_U426_in),
    .clk(_U426_clk),
    .out(_U426_out)
);
assign _U427_in = in[2];
assign _U427_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U427 (
    .in(_U427_in),
    .clk(_U427_clk),
    .out(_U427_out)
);
assign _U428_in = in[3];
assign _U428_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U428_in),
    .clk(_U428_clk),
    .out(_U428_out)
);
assign _U429_in = in[4];
assign _U429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U429 (
    .in(_U429_in),
    .clk(_U429_clk),
    .out(_U429_out)
);
assign out[4] = _U429_out;
assign out[3] = _U428_out;
assign out[2] = _U427_out;
assign out[1] = _U426_out;
assign out[0] = _U425_out;
endmodule

module array_delay_U417 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U418_in;
wire _U418_clk;
wire [15:0] _U418_out;
wire [15:0] _U419_in;
wire _U419_clk;
wire [15:0] _U419_out;
wire [15:0] _U420_in;
wire _U420_clk;
wire [15:0] _U420_out;
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire _U422_clk;
wire [15:0] _U422_out;
assign _U418_in = in[0];
assign _U418_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U418 (
    .in(_U418_in),
    .clk(_U418_clk),
    .out(_U418_out)
);
assign _U419_in = in[1];
assign _U419_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U419 (
    .in(_U419_in),
    .clk(_U419_clk),
    .out(_U419_out)
);
assign _U420_in = in[2];
assign _U420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U420_in),
    .clk(_U420_clk),
    .out(_U420_out)
);
assign _U421_in = in[3];
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = in[4];
assign _U422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U422 (
    .in(_U422_in),
    .clk(_U422_clk),
    .out(_U422_out)
);
assign out[4] = _U422_out;
assign out[3] = _U421_out;
assign out[2] = _U420_out;
assign out[1] = _U419_out;
assign out[0] = _U418_out;
endmodule

module array_delay_U410 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U411_in;
wire _U411_clk;
wire [15:0] _U411_out;
wire [15:0] _U412_in;
wire _U412_clk;
wire [15:0] _U412_out;
wire [15:0] _U413_in;
wire _U413_clk;
wire [15:0] _U413_out;
wire [15:0] _U414_in;
wire _U414_clk;
wire [15:0] _U414_out;
wire [15:0] _U415_in;
wire _U415_clk;
wire [15:0] _U415_out;
assign _U411_in = in[0];
assign _U411_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U411 (
    .in(_U411_in),
    .clk(_U411_clk),
    .out(_U411_out)
);
assign _U412_in = in[1];
assign _U412_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U412 (
    .in(_U412_in),
    .clk(_U412_clk),
    .out(_U412_out)
);
assign _U413_in = in[2];
assign _U413_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U413 (
    .in(_U413_in),
    .clk(_U413_clk),
    .out(_U413_out)
);
assign _U414_in = in[3];
assign _U414_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U414 (
    .in(_U414_in),
    .clk(_U414_clk),
    .out(_U414_out)
);
assign _U415_in = in[4];
assign _U415_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U415 (
    .in(_U415_in),
    .clk(_U415_clk),
    .out(_U415_out)
);
assign out[4] = _U415_out;
assign out[3] = _U414_out;
assign out[2] = _U413_out;
assign out[1] = _U412_out;
assign out[0] = _U411_out;
endmodule

module array_delay_U403 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U404_in;
wire _U404_clk;
wire [15:0] _U404_out;
wire [15:0] _U405_in;
wire _U405_clk;
wire [15:0] _U405_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire _U407_clk;
wire [15:0] _U407_out;
wire [15:0] _U408_in;
wire _U408_clk;
wire [15:0] _U408_out;
assign _U404_in = in[0];
assign _U404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U404 (
    .in(_U404_in),
    .clk(_U404_clk),
    .out(_U404_out)
);
assign _U405_in = in[1];
assign _U405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(_U405_in),
    .clk(_U405_clk),
    .out(_U405_out)
);
assign _U406_in = in[2];
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = in[3];
assign _U407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U407 (
    .in(_U407_in),
    .clk(_U407_clk),
    .out(_U407_out)
);
assign _U408_in = in[4];
assign _U408_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U408 (
    .in(_U408_in),
    .clk(_U408_clk),
    .out(_U408_out)
);
assign out[4] = _U408_out;
assign out[3] = _U407_out;
assign out[2] = _U406_out;
assign out[1] = _U405_out;
assign out[0] = _U404_out;
endmodule

module array_delay_U396 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U397_in;
wire _U397_clk;
wire [15:0] _U397_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
wire [15:0] _U400_in;
wire _U400_clk;
wire [15:0] _U400_out;
wire [15:0] _U401_in;
wire _U401_clk;
wire [15:0] _U401_out;
assign _U397_in = in[0];
assign _U397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U397_in),
    .clk(_U397_clk),
    .out(_U397_out)
);
assign _U398_in = in[1];
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = in[2];
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign _U400_in = in[3];
assign _U400_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U400 (
    .in(_U400_in),
    .clk(_U400_clk),
    .out(_U400_out)
);
assign _U401_in = in[4];
assign _U401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U401_in),
    .clk(_U401_clk),
    .out(_U401_out)
);
assign out[4] = _U401_out;
assign out[3] = _U400_out;
assign out[2] = _U399_out;
assign out[1] = _U398_out;
assign out[0] = _U397_out;
endmodule

module array_delay_U389 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U390_in;
wire _U390_clk;
wire [15:0] _U390_out;
wire [15:0] _U391_in;
wire _U391_clk;
wire [15:0] _U391_out;
wire [15:0] _U392_in;
wire _U392_clk;
wire [15:0] _U392_out;
wire [15:0] _U393_in;
wire _U393_clk;
wire [15:0] _U393_out;
wire [15:0] _U394_in;
wire _U394_clk;
wire [15:0] _U394_out;
assign _U390_in = in[0];
assign _U390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(_U390_in),
    .clk(_U390_clk),
    .out(_U390_out)
);
assign _U391_in = in[1];
assign _U391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U391_in),
    .clk(_U391_clk),
    .out(_U391_out)
);
assign _U392_in = in[2];
assign _U392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U392_in),
    .clk(_U392_clk),
    .out(_U392_out)
);
assign _U393_in = in[3];
assign _U393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U393 (
    .in(_U393_in),
    .clk(_U393_clk),
    .out(_U393_out)
);
assign _U394_in = in[4];
assign _U394_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U394 (
    .in(_U394_in),
    .clk(_U394_clk),
    .out(_U394_out)
);
assign out[4] = _U394_out;
assign out[3] = _U393_out;
assign out[2] = _U392_out;
assign out[1] = _U391_out;
assign out[0] = _U390_out;
endmodule

module array_delay_U382 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U383_in;
wire _U383_clk;
wire [15:0] _U383_out;
wire [15:0] _U384_in;
wire _U384_clk;
wire [15:0] _U384_out;
wire [15:0] _U385_in;
wire _U385_clk;
wire [15:0] _U385_out;
wire [15:0] _U386_in;
wire _U386_clk;
wire [15:0] _U386_out;
wire [15:0] _U387_in;
wire _U387_clk;
wire [15:0] _U387_out;
assign _U383_in = in[0];
assign _U383_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U383 (
    .in(_U383_in),
    .clk(_U383_clk),
    .out(_U383_out)
);
assign _U384_in = in[1];
assign _U384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U384 (
    .in(_U384_in),
    .clk(_U384_clk),
    .out(_U384_out)
);
assign _U385_in = in[2];
assign _U385_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U385 (
    .in(_U385_in),
    .clk(_U385_clk),
    .out(_U385_out)
);
assign _U386_in = in[3];
assign _U386_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U386 (
    .in(_U386_in),
    .clk(_U386_clk),
    .out(_U386_out)
);
assign _U387_in = in[4];
assign _U387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U387 (
    .in(_U387_in),
    .clk(_U387_clk),
    .out(_U387_out)
);
assign out[4] = _U387_out;
assign out[3] = _U386_out;
assign out[2] = _U385_out;
assign out[1] = _U384_out;
assign out[0] = _U383_out;
endmodule

module array_delay_U375 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U376_in;
wire _U376_clk;
wire [15:0] _U376_out;
wire [15:0] _U377_in;
wire _U377_clk;
wire [15:0] _U377_out;
wire [15:0] _U378_in;
wire _U378_clk;
wire [15:0] _U378_out;
wire [15:0] _U379_in;
wire _U379_clk;
wire [15:0] _U379_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
assign _U376_in = in[0];
assign _U376_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U376 (
    .in(_U376_in),
    .clk(_U376_clk),
    .out(_U376_out)
);
assign _U377_in = in[1];
assign _U377_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U377 (
    .in(_U377_in),
    .clk(_U377_clk),
    .out(_U377_out)
);
assign _U378_in = in[2];
assign _U378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U378_in),
    .clk(_U378_clk),
    .out(_U378_out)
);
assign _U379_in = in[3];
assign _U379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U379_in),
    .clk(_U379_clk),
    .out(_U379_out)
);
assign _U380_in = in[4];
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign out[4] = _U380_out;
assign out[3] = _U379_out;
assign out[2] = _U378_out;
assign out[1] = _U377_out;
assign out[0] = _U376_out;
endmodule

module array_delay_U368 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U369_in;
wire _U369_clk;
wire [15:0] _U369_out;
wire [15:0] _U370_in;
wire _U370_clk;
wire [15:0] _U370_out;
wire [15:0] _U371_in;
wire _U371_clk;
wire [15:0] _U371_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire _U373_clk;
wire [15:0] _U373_out;
assign _U369_in = in[0];
assign _U369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U369 (
    .in(_U369_in),
    .clk(_U369_clk),
    .out(_U369_out)
);
assign _U370_in = in[1];
assign _U370_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U370 (
    .in(_U370_in),
    .clk(_U370_clk),
    .out(_U370_out)
);
assign _U371_in = in[2];
assign _U371_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(_U371_in),
    .clk(_U371_clk),
    .out(_U371_out)
);
assign _U372_in = in[3];
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = in[4];
assign _U373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U373 (
    .in(_U373_in),
    .clk(_U373_clk),
    .out(_U373_out)
);
assign out[4] = _U373_out;
assign out[3] = _U372_out;
assign out[2] = _U371_out;
assign out[1] = _U370_out;
assign out[0] = _U369_out;
endmodule

module array_delay_U361 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U362_in;
wire _U362_clk;
wire [15:0] _U362_out;
wire [15:0] _U363_in;
wire _U363_clk;
wire [15:0] _U363_out;
wire [15:0] _U364_in;
wire _U364_clk;
wire [15:0] _U364_out;
wire [15:0] _U365_in;
wire _U365_clk;
wire [15:0] _U365_out;
wire [15:0] _U366_in;
wire _U366_clk;
wire [15:0] _U366_out;
assign _U362_in = in[0];
assign _U362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U362 (
    .in(_U362_in),
    .clk(_U362_clk),
    .out(_U362_out)
);
assign _U363_in = in[1];
assign _U363_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U363 (
    .in(_U363_in),
    .clk(_U363_clk),
    .out(_U363_out)
);
assign _U364_in = in[2];
assign _U364_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U364 (
    .in(_U364_in),
    .clk(_U364_clk),
    .out(_U364_out)
);
assign _U365_in = in[3];
assign _U365_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U365 (
    .in(_U365_in),
    .clk(_U365_clk),
    .out(_U365_out)
);
assign _U366_in = in[4];
assign _U366_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U366 (
    .in(_U366_in),
    .clk(_U366_clk),
    .out(_U366_out)
);
assign out[4] = _U366_out;
assign out[3] = _U365_out;
assign out[2] = _U364_out;
assign out[1] = _U363_out;
assign out[0] = _U362_out;
endmodule

module array_delay_U354 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire _U356_clk;
wire [15:0] _U356_out;
wire [15:0] _U357_in;
wire _U357_clk;
wire [15:0] _U357_out;
wire [15:0] _U358_in;
wire _U358_clk;
wire [15:0] _U358_out;
wire [15:0] _U359_in;
wire _U359_clk;
wire [15:0] _U359_out;
assign _U355_in = in[0];
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = in[1];
assign _U356_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U356 (
    .in(_U356_in),
    .clk(_U356_clk),
    .out(_U356_out)
);
assign _U357_in = in[2];
assign _U357_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U357 (
    .in(_U357_in),
    .clk(_U357_clk),
    .out(_U357_out)
);
assign _U358_in = in[3];
assign _U358_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U358 (
    .in(_U358_in),
    .clk(_U358_clk),
    .out(_U358_out)
);
assign _U359_in = in[4];
assign _U359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U359 (
    .in(_U359_in),
    .clk(_U359_clk),
    .out(_U359_out)
);
assign out[4] = _U359_out;
assign out[3] = _U358_out;
assign out[2] = _U357_out;
assign out[1] = _U356_out;
assign out[0] = _U355_out;
endmodule

module array_delay_U347 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U348_in;
wire _U348_clk;
wire [15:0] _U348_out;
wire [15:0] _U349_in;
wire _U349_clk;
wire [15:0] _U349_out;
wire [15:0] _U350_in;
wire _U350_clk;
wire [15:0] _U350_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire _U352_clk;
wire [15:0] _U352_out;
assign _U348_in = in[0];
assign _U348_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U348 (
    .in(_U348_in),
    .clk(_U348_clk),
    .out(_U348_out)
);
assign _U349_in = in[1];
assign _U349_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U349 (
    .in(_U349_in),
    .clk(_U349_clk),
    .out(_U349_out)
);
assign _U350_in = in[2];
assign _U350_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U350_in),
    .clk(_U350_clk),
    .out(_U350_out)
);
assign _U351_in = in[3];
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = in[4];
assign _U352_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U352 (
    .in(_U352_in),
    .clk(_U352_clk),
    .out(_U352_out)
);
assign out[4] = _U352_out;
assign out[3] = _U351_out;
assign out[2] = _U350_out;
assign out[1] = _U349_out;
assign out[0] = _U348_out;
endmodule

module array_delay_U340 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire _U342_clk;
wire [15:0] _U342_out;
wire [15:0] _U343_in;
wire _U343_clk;
wire [15:0] _U343_out;
wire [15:0] _U344_in;
wire _U344_clk;
wire [15:0] _U344_out;
wire [15:0] _U345_in;
wire _U345_clk;
wire [15:0] _U345_out;
assign _U341_in = in[0];
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = in[1];
assign _U342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U342_in),
    .clk(_U342_clk),
    .out(_U342_out)
);
assign _U343_in = in[2];
assign _U343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U343 (
    .in(_U343_in),
    .clk(_U343_clk),
    .out(_U343_out)
);
assign _U344_in = in[3];
assign _U344_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U344 (
    .in(_U344_in),
    .clk(_U344_clk),
    .out(_U344_out)
);
assign _U345_in = in[4];
assign _U345_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(_U345_in),
    .clk(_U345_clk),
    .out(_U345_out)
);
assign out[4] = _U345_out;
assign out[3] = _U344_out;
assign out[2] = _U343_out;
assign out[1] = _U342_out;
assign out[0] = _U341_out;
endmodule

module array_delay_U333 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U334_in;
wire _U334_clk;
wire [15:0] _U334_out;
wire [15:0] _U335_in;
wire _U335_clk;
wire [15:0] _U335_out;
wire [15:0] _U336_in;
wire _U336_clk;
wire [15:0] _U336_out;
wire [15:0] _U337_in;
wire _U337_clk;
wire [15:0] _U337_out;
wire [15:0] _U338_in;
wire _U338_clk;
wire [15:0] _U338_out;
assign _U334_in = in[0];
assign _U334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U334 (
    .in(_U334_in),
    .clk(_U334_clk),
    .out(_U334_out)
);
assign _U335_in = in[1];
assign _U335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U335 (
    .in(_U335_in),
    .clk(_U335_clk),
    .out(_U335_out)
);
assign _U336_in = in[2];
assign _U336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(_U336_in),
    .clk(_U336_clk),
    .out(_U336_out)
);
assign _U337_in = in[3];
assign _U337_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U337 (
    .in(_U337_in),
    .clk(_U337_clk),
    .out(_U337_out)
);
assign _U338_in = in[4];
assign _U338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U338_in),
    .clk(_U338_clk),
    .out(_U338_out)
);
assign out[4] = _U338_out;
assign out[3] = _U337_out;
assign out[2] = _U336_out;
assign out[1] = _U335_out;
assign out[0] = _U334_out;
endmodule

module array_delay_U307 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire _U310_clk;
wire [15:0] _U310_out;
wire [15:0] _U311_in;
wire _U311_clk;
wire [15:0] _U311_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
assign _U308_in = in[0];
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = in[1];
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = in[2];
assign _U310_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U310 (
    .in(_U310_in),
    .clk(_U310_clk),
    .out(_U310_out)
);
assign _U311_in = in[3];
assign _U311_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U311 (
    .in(_U311_in),
    .clk(_U311_clk),
    .out(_U311_out)
);
assign _U312_in = in[4];
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign out[4] = _U312_out;
assign out[3] = _U311_out;
assign out[2] = _U310_out;
assign out[1] = _U309_out;
assign out[0] = _U308_out;
endmodule

module array_delay_U300 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire _U303_clk;
wire [15:0] _U303_out;
wire [15:0] _U304_in;
wire _U304_clk;
wire [15:0] _U304_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
assign _U301_in = in[0];
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = in[1];
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = in[2];
assign _U303_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U303 (
    .in(_U303_in),
    .clk(_U303_clk),
    .out(_U303_out)
);
assign _U304_in = in[3];
assign _U304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U304 (
    .in(_U304_in),
    .clk(_U304_clk),
    .out(_U304_out)
);
assign _U305_in = in[4];
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign out[4] = _U305_out;
assign out[3] = _U304_out;
assign out[2] = _U303_out;
assign out[1] = _U302_out;
assign out[0] = _U301_out;
endmodule

module array_delay_U234 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U235_in;
wire _U235_clk;
wire [15:0] _U235_out;
wire [15:0] _U236_in;
wire _U236_clk;
wire [15:0] _U236_out;
wire [15:0] _U237_in;
wire _U237_clk;
wire [15:0] _U237_out;
wire [15:0] _U238_in;
wire _U238_clk;
wire [15:0] _U238_out;
wire [15:0] _U239_in;
wire _U239_clk;
wire [15:0] _U239_out;
assign _U235_in = in[0];
assign _U235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U235 (
    .in(_U235_in),
    .clk(_U235_clk),
    .out(_U235_out)
);
assign _U236_in = in[1];
assign _U236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U236 (
    .in(_U236_in),
    .clk(_U236_clk),
    .out(_U236_out)
);
assign _U237_in = in[2];
assign _U237_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U237 (
    .in(_U237_in),
    .clk(_U237_clk),
    .out(_U237_out)
);
assign _U238_in = in[3];
assign _U238_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U238 (
    .in(_U238_in),
    .clk(_U238_clk),
    .out(_U238_out)
);
assign _U239_in = in[4];
assign _U239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U239 (
    .in(_U239_in),
    .clk(_U239_clk),
    .out(_U239_out)
);
assign out[4] = _U239_out;
assign out[3] = _U238_out;
assign out[2] = _U237_out;
assign out[1] = _U236_out;
assign out[0] = _U235_out;
endmodule

module array_delay_U227 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
wire [15:0] _U229_in;
wire _U229_clk;
wire [15:0] _U229_out;
wire [15:0] _U230_in;
wire _U230_clk;
wire [15:0] _U230_out;
wire [15:0] _U231_in;
wire _U231_clk;
wire [15:0] _U231_out;
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
assign _U228_in = in[0];
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign _U229_in = in[1];
assign _U229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U229_in),
    .clk(_U229_clk),
    .out(_U229_out)
);
assign _U230_in = in[2];
assign _U230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U230 (
    .in(_U230_in),
    .clk(_U230_clk),
    .out(_U230_out)
);
assign _U231_in = in[3];
assign _U231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U231 (
    .in(_U231_in),
    .clk(_U231_clk),
    .out(_U231_out)
);
assign _U232_in = in[4];
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign out[4] = _U232_out;
assign out[3] = _U231_out;
assign out[2] = _U230_out;
assign out[1] = _U229_out;
assign out[0] = _U228_out;
endmodule

module array_delay_U220 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
wire [15:0] _U223_in;
wire _U223_clk;
wire [15:0] _U223_out;
wire [15:0] _U224_in;
wire _U224_clk;
wire [15:0] _U224_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
assign _U221_in = in[0];
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign _U222_in = in[1];
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign _U223_in = in[2];
assign _U223_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(_U223_in),
    .clk(_U223_clk),
    .out(_U223_out)
);
assign _U224_in = in[3];
assign _U224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U224_in),
    .clk(_U224_clk),
    .out(_U224_out)
);
assign _U225_in = in[4];
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign out[4] = _U225_out;
assign out[3] = _U224_out;
assign out[2] = _U223_out;
assign out[1] = _U222_out;
assign out[0] = _U221_out;
endmodule

module array_delay_U213 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire _U215_clk;
wire [15:0] _U215_out;
wire [15:0] _U216_in;
wire _U216_clk;
wire [15:0] _U216_out;
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
assign _U214_in = in[0];
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = in[1];
assign _U215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(_U215_in),
    .clk(_U215_clk),
    .out(_U215_out)
);
assign _U216_in = in[2];
assign _U216_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(_U216_in),
    .clk(_U216_clk),
    .out(_U216_out)
);
assign _U217_in = in[3];
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = in[4];
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign out[4] = _U218_out;
assign out[3] = _U217_out;
assign out[2] = _U216_out;
assign out[1] = _U215_out;
assign out[0] = _U214_out;
endmodule

module array_delay_U206 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U207_in;
wire _U207_clk;
wire [15:0] _U207_out;
wire [15:0] _U208_in;
wire _U208_clk;
wire [15:0] _U208_out;
wire [15:0] _U209_in;
wire _U209_clk;
wire [15:0] _U209_out;
wire [15:0] _U210_in;
wire _U210_clk;
wire [15:0] _U210_out;
wire [15:0] _U211_in;
wire _U211_clk;
wire [15:0] _U211_out;
assign _U207_in = in[0];
assign _U207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(_U207_in),
    .clk(_U207_clk),
    .out(_U207_out)
);
assign _U208_in = in[1];
assign _U208_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U208 (
    .in(_U208_in),
    .clk(_U208_clk),
    .out(_U208_out)
);
assign _U209_in = in[2];
assign _U209_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U209 (
    .in(_U209_in),
    .clk(_U209_clk),
    .out(_U209_out)
);
assign _U210_in = in[3];
assign _U210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U210 (
    .in(_U210_in),
    .clk(_U210_clk),
    .out(_U210_out)
);
assign _U211_in = in[4];
assign _U211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(_U211_in),
    .clk(_U211_clk),
    .out(_U211_out)
);
assign out[4] = _U211_out;
assign out[3] = _U210_out;
assign out[2] = _U209_out;
assign out[1] = _U208_out;
assign out[0] = _U207_out;
endmodule

module array_delay_U199 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U200_in;
wire _U200_clk;
wire [15:0] _U200_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
wire [15:0] _U202_in;
wire _U202_clk;
wire [15:0] _U202_out;
wire [15:0] _U203_in;
wire _U203_clk;
wire [15:0] _U203_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
assign _U200_in = in[0];
assign _U200_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U200 (
    .in(_U200_in),
    .clk(_U200_clk),
    .out(_U200_out)
);
assign _U201_in = in[1];
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign _U202_in = in[2];
assign _U202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U202 (
    .in(_U202_in),
    .clk(_U202_clk),
    .out(_U202_out)
);
assign _U203_in = in[3];
assign _U203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U203 (
    .in(_U203_in),
    .clk(_U203_clk),
    .out(_U203_out)
);
assign _U204_in = in[4];
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign out[4] = _U204_out;
assign out[3] = _U203_out;
assign out[2] = _U202_out;
assign out[1] = _U201_out;
assign out[0] = _U200_out;
endmodule

module array_delay_U192 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U193_in;
wire _U193_clk;
wire [15:0] _U193_out;
wire [15:0] _U194_in;
wire _U194_clk;
wire [15:0] _U194_out;
wire [15:0] _U195_in;
wire _U195_clk;
wire [15:0] _U195_out;
wire [15:0] _U196_in;
wire _U196_clk;
wire [15:0] _U196_out;
wire [15:0] _U197_in;
wire _U197_clk;
wire [15:0] _U197_out;
assign _U193_in = in[0];
assign _U193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U193_in),
    .clk(_U193_clk),
    .out(_U193_out)
);
assign _U194_in = in[1];
assign _U194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U194 (
    .in(_U194_in),
    .clk(_U194_clk),
    .out(_U194_out)
);
assign _U195_in = in[2];
assign _U195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U195 (
    .in(_U195_in),
    .clk(_U195_clk),
    .out(_U195_out)
);
assign _U196_in = in[3];
assign _U196_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U196 (
    .in(_U196_in),
    .clk(_U196_clk),
    .out(_U196_out)
);
assign _U197_in = in[4];
assign _U197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U197 (
    .in(_U197_in),
    .clk(_U197_clk),
    .out(_U197_out)
);
assign out[4] = _U197_out;
assign out[3] = _U196_out;
assign out[2] = _U195_out;
assign out[1] = _U194_out;
assign out[0] = _U193_out;
endmodule

module array_delay_U185 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U186_in;
wire _U186_clk;
wire [15:0] _U186_out;
wire [15:0] _U187_in;
wire _U187_clk;
wire [15:0] _U187_out;
wire [15:0] _U188_in;
wire _U188_clk;
wire [15:0] _U188_out;
wire [15:0] _U189_in;
wire _U189_clk;
wire [15:0] _U189_out;
wire [15:0] _U190_in;
wire _U190_clk;
wire [15:0] _U190_out;
assign _U186_in = in[0];
assign _U186_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U186 (
    .in(_U186_in),
    .clk(_U186_clk),
    .out(_U186_out)
);
assign _U187_in = in[1];
assign _U187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U187 (
    .in(_U187_in),
    .clk(_U187_clk),
    .out(_U187_out)
);
assign _U188_in = in[2];
assign _U188_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U188 (
    .in(_U188_in),
    .clk(_U188_clk),
    .out(_U188_out)
);
assign _U189_in = in[3];
assign _U189_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U189 (
    .in(_U189_in),
    .clk(_U189_clk),
    .out(_U189_out)
);
assign _U190_in = in[4];
assign _U190_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U190 (
    .in(_U190_in),
    .clk(_U190_clk),
    .out(_U190_out)
);
assign out[4] = _U190_out;
assign out[3] = _U189_out;
assign out[2] = _U188_out;
assign out[1] = _U187_out;
assign out[0] = _U186_out;
endmodule

module array_delay_U178 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
wire [15:0] _U180_in;
wire _U180_clk;
wire [15:0] _U180_out;
wire [15:0] _U181_in;
wire _U181_clk;
wire [15:0] _U181_out;
wire [15:0] _U182_in;
wire _U182_clk;
wire [15:0] _U182_out;
wire [15:0] _U183_in;
wire _U183_clk;
wire [15:0] _U183_out;
assign _U179_in = in[0];
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign _U180_in = in[1];
assign _U180_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U180 (
    .in(_U180_in),
    .clk(_U180_clk),
    .out(_U180_out)
);
assign _U181_in = in[2];
assign _U181_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U181 (
    .in(_U181_in),
    .clk(_U181_clk),
    .out(_U181_out)
);
assign _U182_in = in[3];
assign _U182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U182_in),
    .clk(_U182_clk),
    .out(_U182_out)
);
assign _U183_in = in[4];
assign _U183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U183_in),
    .clk(_U183_clk),
    .out(_U183_out)
);
assign out[4] = _U183_out;
assign out[3] = _U182_out;
assign out[2] = _U181_out;
assign out[1] = _U180_out;
assign out[0] = _U179_out;
endmodule

module array_delay_U171 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U172_in;
wire _U172_clk;
wire [15:0] _U172_out;
wire [15:0] _U173_in;
wire _U173_clk;
wire [15:0] _U173_out;
wire [15:0] _U174_in;
wire _U174_clk;
wire [15:0] _U174_out;
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
wire [15:0] _U176_in;
wire _U176_clk;
wire [15:0] _U176_out;
assign _U172_in = in[0];
assign _U172_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(_U172_in),
    .clk(_U172_clk),
    .out(_U172_out)
);
assign _U173_in = in[1];
assign _U173_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U173 (
    .in(_U173_in),
    .clk(_U173_clk),
    .out(_U173_out)
);
assign _U174_in = in[2];
assign _U174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(_U174_in),
    .clk(_U174_clk),
    .out(_U174_out)
);
assign _U175_in = in[3];
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign _U176_in = in[4];
assign _U176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U176 (
    .in(_U176_in),
    .clk(_U176_clk),
    .out(_U176_out)
);
assign out[4] = _U176_out;
assign out[3] = _U175_out;
assign out[2] = _U174_out;
assign out[1] = _U173_out;
assign out[0] = _U172_out;
endmodule

module array_delay_U164 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U165_in;
wire _U165_clk;
wire [15:0] _U165_out;
wire [15:0] _U166_in;
wire _U166_clk;
wire [15:0] _U166_out;
wire [15:0] _U167_in;
wire _U167_clk;
wire [15:0] _U167_out;
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
wire [15:0] _U169_in;
wire _U169_clk;
wire [15:0] _U169_out;
assign _U165_in = in[0];
assign _U165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(_U165_in),
    .clk(_U165_clk),
    .out(_U165_out)
);
assign _U166_in = in[1];
assign _U166_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(_U166_in),
    .clk(_U166_clk),
    .out(_U166_out)
);
assign _U167_in = in[2];
assign _U167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U167_in),
    .clk(_U167_clk),
    .out(_U167_out)
);
assign _U168_in = in[3];
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign _U169_in = in[4];
assign _U169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U169 (
    .in(_U169_in),
    .clk(_U169_clk),
    .out(_U169_out)
);
assign out[4] = _U169_out;
assign out[3] = _U168_out;
assign out[2] = _U167_out;
assign out[1] = _U166_out;
assign out[0] = _U165_out;
endmodule

module array_delay_U157 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U158_in;
wire _U158_clk;
wire [15:0] _U158_out;
wire [15:0] _U159_in;
wire _U159_clk;
wire [15:0] _U159_out;
wire [15:0] _U160_in;
wire _U160_clk;
wire [15:0] _U160_out;
wire [15:0] _U161_in;
wire _U161_clk;
wire [15:0] _U161_out;
wire [15:0] _U162_in;
wire _U162_clk;
wire [15:0] _U162_out;
assign _U158_in = in[0];
assign _U158_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U158 (
    .in(_U158_in),
    .clk(_U158_clk),
    .out(_U158_out)
);
assign _U159_in = in[1];
assign _U159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U159_in),
    .clk(_U159_clk),
    .out(_U159_out)
);
assign _U160_in = in[2];
assign _U160_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U160 (
    .in(_U160_in),
    .clk(_U160_clk),
    .out(_U160_out)
);
assign _U161_in = in[3];
assign _U161_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U161 (
    .in(_U161_in),
    .clk(_U161_clk),
    .out(_U161_out)
);
assign _U162_in = in[4];
assign _U162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(_U162_in),
    .clk(_U162_clk),
    .out(_U162_out)
);
assign out[4] = _U162_out;
assign out[3] = _U161_out;
assign out[2] = _U160_out;
assign out[1] = _U159_out;
assign out[0] = _U158_out;
endmodule

module array_delay_U150 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U151_in;
wire _U151_clk;
wire [15:0] _U151_out;
wire [15:0] _U152_in;
wire _U152_clk;
wire [15:0] _U152_out;
wire [15:0] _U153_in;
wire _U153_clk;
wire [15:0] _U153_out;
wire [15:0] _U154_in;
wire _U154_clk;
wire [15:0] _U154_out;
wire [15:0] _U155_in;
wire _U155_clk;
wire [15:0] _U155_out;
assign _U151_in = in[0];
assign _U151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(_U151_in),
    .clk(_U151_clk),
    .out(_U151_out)
);
assign _U152_in = in[1];
assign _U152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U152 (
    .in(_U152_in),
    .clk(_U152_clk),
    .out(_U152_out)
);
assign _U153_in = in[2];
assign _U153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U153 (
    .in(_U153_in),
    .clk(_U153_clk),
    .out(_U153_out)
);
assign _U154_in = in[3];
assign _U154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(_U154_in),
    .clk(_U154_clk),
    .out(_U154_out)
);
assign _U155_in = in[4];
assign _U155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U155_in),
    .clk(_U155_clk),
    .out(_U155_out)
);
assign out[4] = _U155_out;
assign out[3] = _U154_out;
assign out[2] = _U153_out;
assign out[1] = _U152_out;
assign out[0] = _U151_out;
endmodule

module array_delay_U143 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U144_in;
wire _U144_clk;
wire [15:0] _U144_out;
wire [15:0] _U145_in;
wire _U145_clk;
wire [15:0] _U145_out;
wire [15:0] _U146_in;
wire _U146_clk;
wire [15:0] _U146_out;
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire _U148_clk;
wire [15:0] _U148_out;
assign _U144_in = in[0];
assign _U144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U144 (
    .in(_U144_in),
    .clk(_U144_clk),
    .out(_U144_out)
);
assign _U145_in = in[1];
assign _U145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U145_in),
    .clk(_U145_clk),
    .out(_U145_out)
);
assign _U146_in = in[2];
assign _U146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U146_in),
    .clk(_U146_clk),
    .out(_U146_out)
);
assign _U147_in = in[3];
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = in[4];
assign _U148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U148_in),
    .clk(_U148_clk),
    .out(_U148_out)
);
assign out[4] = _U148_out;
assign out[3] = _U147_out;
assign out[2] = _U146_out;
assign out[1] = _U145_out;
assign out[0] = _U144_out;
endmodule

module array_delay_U136 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U137_in;
wire _U137_clk;
wire [15:0] _U137_out;
wire [15:0] _U138_in;
wire _U138_clk;
wire [15:0] _U138_out;
wire [15:0] _U139_in;
wire _U139_clk;
wire [15:0] _U139_out;
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire _U141_clk;
wire [15:0] _U141_out;
assign _U137_in = in[0];
assign _U137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U137 (
    .in(_U137_in),
    .clk(_U137_clk),
    .out(_U137_out)
);
assign _U138_in = in[1];
assign _U138_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U138 (
    .in(_U138_in),
    .clk(_U138_clk),
    .out(_U138_out)
);
assign _U139_in = in[2];
assign _U139_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U139 (
    .in(_U139_in),
    .clk(_U139_clk),
    .out(_U139_out)
);
assign _U140_in = in[3];
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = in[4];
assign _U141_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U141 (
    .in(_U141_in),
    .clk(_U141_clk),
    .out(_U141_out)
);
assign out[4] = _U141_out;
assign out[3] = _U140_out;
assign out[2] = _U139_out;
assign out[1] = _U138_out;
assign out[0] = _U137_out;
endmodule

module array_delay_U129 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U130_in;
wire _U130_clk;
wire [15:0] _U130_out;
wire [15:0] _U131_in;
wire _U131_clk;
wire [15:0] _U131_out;
wire [15:0] _U132_in;
wire _U132_clk;
wire [15:0] _U132_out;
wire [15:0] _U133_in;
wire _U133_clk;
wire [15:0] _U133_out;
wire [15:0] _U134_in;
wire _U134_clk;
wire [15:0] _U134_out;
assign _U130_in = in[0];
assign _U130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U130_in),
    .clk(_U130_clk),
    .out(_U130_out)
);
assign _U131_in = in[1];
assign _U131_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U131 (
    .in(_U131_in),
    .clk(_U131_clk),
    .out(_U131_out)
);
assign _U132_in = in[2];
assign _U132_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(_U132_in),
    .clk(_U132_clk),
    .out(_U132_out)
);
assign _U133_in = in[3];
assign _U133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U133_in),
    .clk(_U133_clk),
    .out(_U133_out)
);
assign _U134_in = in[4];
assign _U134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U134_in),
    .clk(_U134_clk),
    .out(_U134_out)
);
assign out[4] = _U134_out;
assign out[3] = _U133_out;
assign out[2] = _U132_out;
assign out[1] = _U131_out;
assign out[0] = _U130_out;
endmodule

module array_delay_U122 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
wire [15:0] _U125_in;
wire _U125_clk;
wire [15:0] _U125_out;
wire [15:0] _U126_in;
wire _U126_clk;
wire [15:0] _U126_out;
wire [15:0] _U127_in;
wire _U127_clk;
wire [15:0] _U127_out;
assign _U123_in = in[0];
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = in[1];
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign _U125_in = in[2];
assign _U125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U125 (
    .in(_U125_in),
    .clk(_U125_clk),
    .out(_U125_out)
);
assign _U126_in = in[3];
assign _U126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(_U126_in),
    .clk(_U126_clk),
    .out(_U126_out)
);
assign _U127_in = in[4];
assign _U127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U127_in),
    .clk(_U127_clk),
    .out(_U127_out)
);
assign out[4] = _U127_out;
assign out[3] = _U126_out;
assign out[2] = _U125_out;
assign out[1] = _U124_out;
assign out[0] = _U123_out;
endmodule

module aff__U699 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h032c * d[1])))) + (16'(16'h001d * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h7d21);
endmodule

module affine_controller__U698 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U699 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U663 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0051 * d[1])))) + (16'(16'h001b * d[2])))) + (16'(16'h0009 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U662 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U663 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0002;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U53 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U52 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U53 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U475 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U474 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U475 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U452 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U451 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U452 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U30 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U29 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U30 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U264 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U263 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U264 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U241 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U240 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U241 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h010e * d[1])))) + (16'(16'h0009 * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h0001);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module _U88_pt__U89 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U85_pt__U86 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U81_pt__U82 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U7_pt__U8 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U78_pt__U79 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U72_pt__U73 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U69_pt__U70 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U61_pt__U62 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U613_pt__U614 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U613_in;
assign _U613_in = in0_conv_stencil[0];
_U613_pt__U614 _U613 (
    .in(_U613_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U611_pt__U612 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_kernel_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
wire [15:0] _U611_in;
assign _U611_in = in0_hw_kernel_stencil[0];
_U611_pt__U612 _U611 (
    .in(_U611_in),
    .out(out_hw_kernel_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module _U594_pt__U595 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U58_pt__U59 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U585_pt__U586 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U576_pt__U577 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U568_pt__U569 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U560_pt__U561 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U553_pt__U554 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U546_pt__U547 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U540_pt__U541 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U534_pt__U535 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U529_pt__U530 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U524_pt__U525 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U520_pt__U521 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U516_pt__U517 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U513_pt__U514 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U510_pt__U511 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U508_pt__U509 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U506_pt__U507 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U4_pt__U5 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U490_pt__U491 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U48_pt__U49 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U487_pt__U488 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U483_pt__U484 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U480_pt__U481 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U474_pt__U475 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U471_pt__U472 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U463_pt__U464 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U460_pt__U461 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U45_pt__U46 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U450_pt__U451 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U447_pt__U448 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U435_pt__U436 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U432_pt__U433 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U429_pt__U430 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U415_pt__U416 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U413_pt__U414 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U410_pt__U411 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_3_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U410_in;
wire [15:0] _U410_out;
wire [15:0] _U412_in;
wire _U412_clk;
wire [15:0] _U412_out;
wire [15:0] _U413_in;
wire [15:0] _U415_in;
wire [15:0] _U415_out;
wire [15:0] _U417_in;
wire _U417_clk;
wire [15:0] _U417_out;
wire [15:0] _U418_in;
wire _U418_clk;
wire [15:0] _U418_out;
wire [15:0] _U419_in;
wire _U419_clk;
wire [15:0] _U419_out;
wire [15:0] _U420_in;
wire _U420_clk;
wire [15:0] _U420_out;
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire _U422_clk;
wire [15:0] _U422_out;
wire [15:0] _U423_in;
wire _U423_clk;
wire [15:0] _U423_out;
wire [15:0] _U424_in;
wire _U424_clk;
wire [15:0] _U424_out;
wire [15:0] _U425_in;
wire _U425_clk;
wire [15:0] _U425_out;
wire [15:0] _U426_in;
wire _U426_clk;
wire [15:0] _U426_out;
wire [15:0] _U427_in;
wire _U427_clk;
wire [15:0] _U427_out;
wire [15:0] _U428_in;
wire _U428_clk;
wire [15:0] _U428_out;
wire [15:0] _U429_in;
wire [15:0] _U429_out;
wire [15:0] _U431_in;
wire _U431_clk;
wire [15:0] _U431_out;
wire [15:0] _U432_in;
wire [15:0] _U432_out;
wire [15:0] _U434_in;
wire _U434_clk;
wire [15:0] _U434_out;
wire [15:0] _U435_in;
wire [15:0] _U435_out;
wire [15:0] _U437_in;
wire _U437_clk;
wire [15:0] _U437_out;
wire [15:0] _U438_in;
wire _U438_clk;
wire [15:0] _U438_out;
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
wire [15:0] _U447_in;
wire [15:0] _U447_out;
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire [15:0] _U450_out;
wire [15:0] _U452_in;
wire _U452_clk;
wire [15:0] _U452_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
wire [15:0] _U454_in;
wire _U454_clk;
wire [15:0] _U454_out;
wire [15:0] _U455_in;
wire _U455_clk;
wire [15:0] _U455_out;
wire [15:0] _U456_in;
wire _U456_clk;
wire [15:0] _U456_out;
wire [15:0] _U457_in;
wire _U457_clk;
wire [15:0] _U457_out;
wire [15:0] _U458_in;
wire _U458_clk;
wire [15:0] _U458_out;
wire [15:0] _U459_in;
wire _U459_clk;
wire [15:0] _U459_out;
wire [15:0] _U460_in;
wire [15:0] _U460_out;
wire [15:0] _U462_in;
wire _U462_clk;
wire [15:0] _U462_out;
wire [15:0] _U463_in;
wire [15:0] _U463_out;
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire _U466_clk;
wire [15:0] _U466_out;
wire [15:0] _U467_in;
wire _U467_clk;
wire [15:0] _U467_out;
wire [15:0] _U468_in;
wire _U468_clk;
wire [15:0] _U468_out;
wire [15:0] _U469_in;
wire _U469_clk;
wire [15:0] _U469_out;
wire [15:0] _U470_in;
wire _U470_clk;
wire [15:0] _U470_out;
wire [15:0] _U471_in;
wire [15:0] _U471_out;
wire [15:0] _U473_in;
wire _U473_clk;
wire [15:0] _U473_out;
wire [15:0] _U474_in;
wire [15:0] _U474_out;
wire [15:0] _U476_in;
wire _U476_clk;
wire [15:0] _U476_out;
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire _U478_clk;
wire [15:0] _U478_out;
wire [15:0] _U479_in;
wire _U479_clk;
wire [15:0] _U479_out;
wire [15:0] _U480_in;
wire [15:0] _U480_out;
wire [15:0] _U482_in;
wire _U482_clk;
wire [15:0] _U482_out;
wire [15:0] _U483_in;
wire [15:0] _U483_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire [15:0] _U487_out;
wire [15:0] _U489_in;
wire _U489_clk;
wire [15:0] _U489_out;
wire [15:0] _U490_in;
wire [15:0] _U490_out;
wire [15:0] _U492_in;
wire _U492_clk;
wire [15:0] _U492_out;
wire [15:0] _U493_in;
wire _U493_clk;
wire [15:0] _U493_out;
wire [15:0] _U494_in;
wire _U494_clk;
wire [15:0] _U494_out;
wire [15:0] _U495_in;
wire _U495_clk;
wire [15:0] _U495_out;
wire [15:0] _U496_in;
wire _U496_clk;
wire [15:0] _U496_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
wire [15:0] _U498_in;
wire _U498_clk;
wire [15:0] _U498_out;
wire [15:0] _U499_in;
wire _U499_clk;
wire [15:0] _U499_out;
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire _U502_clk;
wire [15:0] _U502_out;
wire [15:0] _U503_in;
wire _U503_clk;
wire [15:0] _U503_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire [15:0] _U506_out;
wire [15:0] _U508_in;
wire [15:0] _U508_out;
wire [15:0] _U510_in;
wire [15:0] _U510_out;
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire [15:0] _U513_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire [15:0] _U516_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire [15:0] _U520_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
wire [15:0] _U524_in;
wire [15:0] _U524_out;
wire [15:0] _U526_in;
wire _U526_clk;
wire [15:0] _U526_out;
wire [15:0] _U527_in;
wire _U527_clk;
wire [15:0] _U527_out;
wire [15:0] _U528_in;
wire _U528_clk;
wire [15:0] _U528_out;
wire [15:0] _U529_in;
wire [15:0] _U529_out;
wire [15:0] _U531_in;
wire _U531_clk;
wire [15:0] _U531_out;
wire [15:0] _U532_in;
wire _U532_clk;
wire [15:0] _U532_out;
wire [15:0] _U533_in;
wire _U533_clk;
wire [15:0] _U533_out;
wire [15:0] _U534_in;
wire [15:0] _U534_out;
wire [15:0] _U536_in;
wire _U536_clk;
wire [15:0] _U536_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire _U539_clk;
wire [15:0] _U539_out;
wire [15:0] _U540_in;
wire [15:0] _U540_out;
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
wire [15:0] _U543_in;
wire _U543_clk;
wire [15:0] _U543_out;
wire [15:0] _U544_in;
wire _U544_clk;
wire [15:0] _U544_out;
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire [15:0] _U546_out;
wire [15:0] _U548_in;
wire _U548_clk;
wire [15:0] _U548_out;
wire [15:0] _U549_in;
wire _U549_clk;
wire [15:0] _U549_out;
wire [15:0] _U550_in;
wire _U550_clk;
wire [15:0] _U550_out;
wire [15:0] _U551_in;
wire _U551_clk;
wire [15:0] _U551_out;
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire [15:0] _U553_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
wire [15:0] _U557_in;
wire _U557_clk;
wire [15:0] _U557_out;
wire [15:0] _U558_in;
wire _U558_clk;
wire [15:0] _U558_out;
wire [15:0] _U559_in;
wire _U559_clk;
wire [15:0] _U559_out;
wire [15:0] _U560_in;
wire [15:0] _U560_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
wire [15:0] _U564_in;
wire _U564_clk;
wire [15:0] _U564_out;
wire [15:0] _U565_in;
wire _U565_clk;
wire [15:0] _U565_out;
wire [15:0] _U566_in;
wire _U566_clk;
wire [15:0] _U566_out;
wire [15:0] _U567_in;
wire _U567_clk;
wire [15:0] _U567_out;
wire [15:0] _U568_in;
wire [15:0] _U568_out;
wire [15:0] _U570_in;
wire _U570_clk;
wire [15:0] _U570_out;
wire [15:0] _U571_in;
wire _U571_clk;
wire [15:0] _U571_out;
wire [15:0] _U572_in;
wire _U572_clk;
wire [15:0] _U572_out;
wire [15:0] _U573_in;
wire _U573_clk;
wire [15:0] _U573_out;
wire [15:0] _U574_in;
wire _U574_clk;
wire [15:0] _U574_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire [15:0] _U576_out;
wire [15:0] _U578_in;
wire _U578_clk;
wire [15:0] _U578_out;
wire [15:0] _U579_in;
wire _U579_clk;
wire [15:0] _U579_out;
wire [15:0] _U580_in;
wire _U580_clk;
wire [15:0] _U580_out;
wire [15:0] _U581_in;
wire _U581_clk;
wire [15:0] _U581_out;
wire [15:0] _U582_in;
wire _U582_clk;
wire [15:0] _U582_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
wire [15:0] _U585_in;
wire [15:0] _U585_out;
wire [15:0] _U587_in;
wire _U587_clk;
wire [15:0] _U587_out;
wire [15:0] _U588_in;
wire _U588_clk;
wire [15:0] _U588_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
wire [15:0] _U592_in;
wire _U592_clk;
wire [15:0] _U592_out;
wire [15:0] _U593_in;
wire _U593_clk;
wire [15:0] _U593_out;
wire [15:0] _U594_in;
wire [15:0] _U594_out;
wire [15:0] _U596_in;
wire _U596_clk;
wire [15:0] _U596_out;
wire [15:0] _U597_in;
wire _U597_clk;
wire [15:0] _U597_out;
wire [15:0] _U598_in;
wire _U598_clk;
wire [15:0] _U598_out;
wire [15:0] _U599_in;
wire _U599_clk;
wire [15:0] _U599_out;
wire [15:0] _U600_in;
wire _U600_clk;
wire [15:0] _U600_out;
wire [15:0] _U601_in;
wire _U601_clk;
wire [15:0] _U601_out;
wire [15:0] _U602_in;
wire _U602_clk;
wire [15:0] _U602_out;
wire [15:0] _U603_in;
wire _U603_clk;
wire [15:0] _U603_out;
wire [15:0] _U604_in;
wire _U604_clk;
wire [15:0] _U604_out;
wire [15:0] _U605_in;
wire _U605_clk;
wire [15:0] _U605_out;
wire [15:0] _U606_in;
wire _U606_clk;
wire [15:0] _U606_out;
wire [15:0] _U607_in;
wire _U607_clk;
wire [15:0] _U607_out;
wire [15:0] _U608_in;
wire _U608_clk;
wire [15:0] _U608_out;
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
assign _U410_in = _U412_out;
_U410_pt__U411 _U410 (
    .in(_U410_in),
    .out(_U410_out)
);
assign _U412_in = 16'(_U490_out + _U432_out);
assign _U412_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U412 (
    .in(_U412_in),
    .clk(_U412_clk),
    .out(_U412_out)
);
assign _U413_in = 16'(_U594_out + _U410_out);
_U413_pt__U414 _U413 (
    .in(_U413_in),
    .out(out_conv_stencil)
);
assign _U415_in = _U428_out;
_U415_pt__U416 _U415 (
    .in(_U415_in),
    .out(_U415_out)
);
assign _U417_in = 16'(_U510_out * _U513_out);
assign _U417_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U417 (
    .in(_U417_in),
    .clk(_U417_clk),
    .out(_U417_out)
);
assign _U418_in = _U417_out;
assign _U418_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U418 (
    .in(_U418_in),
    .clk(_U418_clk),
    .out(_U418_out)
);
assign _U419_in = _U418_out;
assign _U419_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U419 (
    .in(_U419_in),
    .clk(_U419_clk),
    .out(_U419_out)
);
assign _U420_in = _U419_out;
assign _U420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U420_in),
    .clk(_U420_clk),
    .out(_U420_out)
);
assign _U421_in = _U420_out;
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = _U421_out;
assign _U422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U422 (
    .in(_U422_in),
    .clk(_U422_clk),
    .out(_U422_out)
);
assign _U423_in = _U422_out;
assign _U423_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U423 (
    .in(_U423_in),
    .clk(_U423_clk),
    .out(_U423_out)
);
assign _U424_in = _U423_out;
assign _U424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U424 (
    .in(_U424_in),
    .clk(_U424_clk),
    .out(_U424_out)
);
assign _U425_in = _U424_out;
assign _U425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U425 (
    .in(_U425_in),
    .clk(_U425_clk),
    .out(_U425_out)
);
assign _U426_in = _U425_out;
assign _U426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U426 (
    .in(_U426_in),
    .clk(_U426_clk),
    .out(_U426_out)
);
assign _U427_in = _U426_out;
assign _U427_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U427 (
    .in(_U427_in),
    .clk(_U427_clk),
    .out(_U427_out)
);
assign _U428_in = _U427_out;
assign _U428_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U428_in),
    .clk(_U428_clk),
    .out(_U428_out)
);
assign _U429_in = _U431_out;
_U429_pt__U430 _U429 (
    .in(_U429_in),
    .out(_U429_out)
);
assign _U431_in = 16'(_U435_out + _U447_out);
assign _U431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U431_in),
    .clk(_U431_clk),
    .out(_U431_out)
);
assign _U432_in = _U434_out;
_U432_pt__U433 _U432 (
    .in(_U432_in),
    .out(_U432_out)
);
assign _U434_in = 16'(_U415_out + _U429_out);
assign _U434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U434_in),
    .clk(_U434_clk),
    .out(_U434_out)
);
assign _U435_in = _U446_out;
_U435_pt__U436 _U435 (
    .in(_U435_in),
    .out(_U435_out)
);
assign _U437_in = 16'(_U516_out * _U520_out);
assign _U437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U437 (
    .in(_U437_in),
    .clk(_U437_clk),
    .out(_U437_out)
);
assign _U438_in = _U437_out;
assign _U438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(_U438_in),
    .clk(_U438_clk),
    .out(_U438_out)
);
assign _U439_in = _U438_out;
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign _U440_in = _U439_out;
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = _U440_out;
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign _U442_in = _U441_out;
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = _U442_out;
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = _U443_out;
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = _U444_out;
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = _U445_out;
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign _U447_in = _U449_out;
_U447_pt__U448 _U447 (
    .in(_U447_in),
    .out(_U447_out)
);
assign _U449_in = 16'(_U450_out + _U460_out);
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = _U459_out;
_U450_pt__U451 _U450 (
    .in(_U450_in),
    .out(_U450_out)
);
assign _U452_in = 16'(_U524_out * _U529_out);
assign _U452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U452_in),
    .clk(_U452_clk),
    .out(_U452_out)
);
assign _U453_in = _U452_out;
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign _U454_in = _U453_out;
assign _U454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U454 (
    .in(_U454_in),
    .clk(_U454_clk),
    .out(_U454_out)
);
assign _U455_in = _U454_out;
assign _U455_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U455 (
    .in(_U455_in),
    .clk(_U455_clk),
    .out(_U455_out)
);
assign _U456_in = _U455_out;
assign _U456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U456 (
    .in(_U456_in),
    .clk(_U456_clk),
    .out(_U456_out)
);
assign _U457_in = _U456_out;
assign _U457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U457 (
    .in(_U457_in),
    .clk(_U457_clk),
    .out(_U457_out)
);
assign _U458_in = _U457_out;
assign _U458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U458 (
    .in(_U458_in),
    .clk(_U458_clk),
    .out(_U458_out)
);
assign _U459_in = _U458_out;
assign _U459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U459 (
    .in(_U459_in),
    .clk(_U459_clk),
    .out(_U459_out)
);
assign _U460_in = _U462_out;
_U460_pt__U461 _U460 (
    .in(_U460_in),
    .out(_U460_out)
);
assign _U462_in = 16'(_U463_out + _U471_out);
assign _U462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U462_in),
    .clk(_U462_clk),
    .out(_U462_out)
);
assign _U463_in = _U470_out;
_U463_pt__U464 _U463 (
    .in(_U463_in),
    .out(_U463_out)
);
assign _U465_in = 16'(_U534_out * _U540_out);
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = _U465_out;
assign _U466_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U466 (
    .in(_U466_in),
    .clk(_U466_clk),
    .out(_U466_out)
);
assign _U467_in = _U466_out;
assign _U467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U467 (
    .in(_U467_in),
    .clk(_U467_clk),
    .out(_U467_out)
);
assign _U468_in = _U467_out;
assign _U468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U468_in),
    .clk(_U468_clk),
    .out(_U468_out)
);
assign _U469_in = _U468_out;
assign _U469_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U469 (
    .in(_U469_in),
    .clk(_U469_clk),
    .out(_U469_out)
);
assign _U470_in = _U469_out;
assign _U470_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U470 (
    .in(_U470_in),
    .clk(_U470_clk),
    .out(_U470_out)
);
assign _U471_in = _U473_out;
_U471_pt__U472 _U471 (
    .in(_U471_in),
    .out(_U471_out)
);
assign _U473_in = 16'(_U474_out + _U480_out);
assign _U473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U473 (
    .in(_U473_in),
    .clk(_U473_clk),
    .out(_U473_out)
);
assign _U474_in = _U479_out;
_U474_pt__U475 _U474 (
    .in(_U474_in),
    .out(_U474_out)
);
assign _U476_in = 16'(_U546_out * _U553_out);
assign _U476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(_U476_in),
    .clk(_U476_clk),
    .out(_U476_out)
);
assign _U477_in = _U476_out;
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = _U477_out;
assign _U478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(_U478_in),
    .clk(_U478_clk),
    .out(_U478_out)
);
assign _U479_in = _U478_out;
assign _U479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(_U479_in),
    .clk(_U479_clk),
    .out(_U479_out)
);
assign _U480_in = _U482_out;
_U480_pt__U481 _U480 (
    .in(_U480_in),
    .out(_U480_out)
);
assign _U482_in = 16'(_U483_out + _U487_out);
assign _U482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U482_in),
    .clk(_U482_clk),
    .out(_U482_out)
);
assign _U483_in = _U486_out;
_U483_pt__U484 _U483 (
    .in(_U483_in),
    .out(_U483_out)
);
assign _U485_in = 16'(_U560_out * _U568_out);
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = _U485_out;
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = _U489_out;
_U487_pt__U488 _U487 (
    .in(_U487_in),
    .out(_U487_out)
);
assign _U489_in = 16'(_U576_out * _U585_out);
assign _U489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U489_in),
    .clk(_U489_clk),
    .out(_U489_out)
);
assign _U490_in = _U505_out;
_U490_pt__U491 _U490 (
    .in(_U490_in),
    .out(_U490_out)
);
assign _U492_in = in0_conv_stencil[0];
assign _U492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(_U492_in),
    .clk(_U492_clk),
    .out(_U492_out)
);
assign _U493_in = _U492_out;
assign _U493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U493 (
    .in(_U493_in),
    .clk(_U493_clk),
    .out(_U493_out)
);
assign _U494_in = _U493_out;
assign _U494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U494 (
    .in(_U494_in),
    .clk(_U494_clk),
    .out(_U494_out)
);
assign _U495_in = _U494_out;
assign _U495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U495 (
    .in(_U495_in),
    .clk(_U495_clk),
    .out(_U495_out)
);
assign _U496_in = _U495_out;
assign _U496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(_U496_in),
    .clk(_U496_clk),
    .out(_U496_out)
);
assign _U497_in = _U496_out;
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign _U498_in = _U497_out;
assign _U498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U498_in),
    .clk(_U498_clk),
    .out(_U498_out)
);
assign _U499_in = _U498_out;
assign _U499_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(_U499_in),
    .clk(_U499_clk),
    .out(_U499_out)
);
assign _U500_in = _U499_out;
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign _U501_in = _U500_out;
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = _U501_out;
assign _U502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U502_in),
    .clk(_U502_clk),
    .out(_U502_out)
);
assign _U503_in = _U502_out;
assign _U503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(_U503_in),
    .clk(_U503_clk),
    .out(_U503_out)
);
assign _U504_in = _U503_out;
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign _U505_in = _U504_out;
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = in2_hw_kernel_global_wrapper_stencil[0];
_U506_pt__U507 _U506 (
    .in(_U506_in),
    .out(_U506_out)
);
assign _U508_in = in1_hw_input_global_wrapper_stencil[0];
_U508_pt__U509 _U508 (
    .in(_U508_in),
    .out(_U508_out)
);
assign _U510_in = _U512_out;
_U510_pt__U511 _U510 (
    .in(_U510_in),
    .out(_U510_out)
);
assign _U512_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = _U515_out;
_U513_pt__U514 _U513 (
    .in(_U513_in),
    .out(_U513_out)
);
assign _U515_in = in1_hw_input_global_wrapper_stencil[1];
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = _U519_out;
_U516_pt__U517 _U516 (
    .in(_U516_in),
    .out(_U516_out)
);
assign _U518_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign _U519_in = _U518_out;
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = _U523_out;
_U520_pt__U521 _U520 (
    .in(_U520_in),
    .out(_U520_out)
);
assign _U522_in = in1_hw_input_global_wrapper_stencil[2];
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = _U522_out;
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign _U524_in = _U528_out;
_U524_pt__U525 _U524 (
    .in(_U524_in),
    .out(_U524_out)
);
assign _U526_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(_U526_in),
    .clk(_U526_clk),
    .out(_U526_out)
);
assign _U527_in = _U526_out;
assign _U527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(_U527_in),
    .clk(_U527_clk),
    .out(_U527_out)
);
assign _U528_in = _U527_out;
assign _U528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(_U528_in),
    .clk(_U528_clk),
    .out(_U528_out)
);
assign _U529_in = _U533_out;
_U529_pt__U530 _U529 (
    .in(_U529_in),
    .out(_U529_out)
);
assign _U531_in = in1_hw_input_global_wrapper_stencil[3];
assign _U531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(_U531_in),
    .clk(_U531_clk),
    .out(_U531_out)
);
assign _U532_in = _U531_out;
assign _U532_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(_U532_in),
    .clk(_U532_clk),
    .out(_U532_out)
);
assign _U533_in = _U532_out;
assign _U533_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U533 (
    .in(_U533_in),
    .clk(_U533_clk),
    .out(_U533_out)
);
assign _U534_in = _U539_out;
_U534_pt__U535 _U534 (
    .in(_U534_in),
    .out(_U534_out)
);
assign _U536_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U536_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U536_in),
    .clk(_U536_clk),
    .out(_U536_out)
);
assign _U537_in = _U536_out;
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign _U538_in = _U537_out;
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = _U538_out;
assign _U539_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U539_in),
    .clk(_U539_clk),
    .out(_U539_out)
);
assign _U540_in = _U545_out;
_U540_pt__U541 _U540 (
    .in(_U540_in),
    .out(_U540_out)
);
assign _U542_in = in1_hw_input_global_wrapper_stencil[4];
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign _U543_in = _U542_out;
assign _U543_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U543 (
    .in(_U543_in),
    .clk(_U543_clk),
    .out(_U543_out)
);
assign _U544_in = _U543_out;
assign _U544_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U544 (
    .in(_U544_in),
    .clk(_U544_clk),
    .out(_U544_out)
);
assign _U545_in = _U544_out;
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = _U552_out;
_U546_pt__U547 _U546 (
    .in(_U546_in),
    .out(_U546_out)
);
assign _U548_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U548_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U548 (
    .in(_U548_in),
    .clk(_U548_clk),
    .out(_U548_out)
);
assign _U549_in = _U548_out;
assign _U549_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U549 (
    .in(_U549_in),
    .clk(_U549_clk),
    .out(_U549_out)
);
assign _U550_in = _U549_out;
assign _U550_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U550 (
    .in(_U550_in),
    .clk(_U550_clk),
    .out(_U550_out)
);
assign _U551_in = _U550_out;
assign _U551_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U551 (
    .in(_U551_in),
    .clk(_U551_clk),
    .out(_U551_out)
);
assign _U552_in = _U551_out;
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = _U559_out;
_U553_pt__U554 _U553 (
    .in(_U553_in),
    .out(_U553_out)
);
assign _U555_in = in1_hw_input_global_wrapper_stencil[5];
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = _U555_out;
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign _U557_in = _U556_out;
assign _U557_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U557 (
    .in(_U557_in),
    .clk(_U557_clk),
    .out(_U557_out)
);
assign _U558_in = _U557_out;
assign _U558_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U558 (
    .in(_U558_in),
    .clk(_U558_clk),
    .out(_U558_out)
);
assign _U559_in = _U558_out;
assign _U559_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U559 (
    .in(_U559_in),
    .clk(_U559_clk),
    .out(_U559_out)
);
assign _U560_in = _U567_out;
_U560_pt__U561 _U560 (
    .in(_U560_in),
    .out(_U560_out)
);
assign _U562_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = _U562_out;
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign _U564_in = _U563_out;
assign _U564_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U564 (
    .in(_U564_in),
    .clk(_U564_clk),
    .out(_U564_out)
);
assign _U565_in = _U564_out;
assign _U565_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U565 (
    .in(_U565_in),
    .clk(_U565_clk),
    .out(_U565_out)
);
assign _U566_in = _U565_out;
assign _U566_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U566 (
    .in(_U566_in),
    .clk(_U566_clk),
    .out(_U566_out)
);
assign _U567_in = _U566_out;
assign _U567_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U567 (
    .in(_U567_in),
    .clk(_U567_clk),
    .out(_U567_out)
);
assign _U568_in = _U575_out;
_U568_pt__U569 _U568 (
    .in(_U568_in),
    .out(_U568_out)
);
assign _U570_in = in1_hw_input_global_wrapper_stencil[6];
assign _U570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U570_in),
    .clk(_U570_clk),
    .out(_U570_out)
);
assign _U571_in = _U570_out;
assign _U571_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U571 (
    .in(_U571_in),
    .clk(_U571_clk),
    .out(_U571_out)
);
assign _U572_in = _U571_out;
assign _U572_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U572 (
    .in(_U572_in),
    .clk(_U572_clk),
    .out(_U572_out)
);
assign _U573_in = _U572_out;
assign _U573_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U573 (
    .in(_U573_in),
    .clk(_U573_clk),
    .out(_U573_out)
);
assign _U574_in = _U573_out;
assign _U574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(_U574_in),
    .clk(_U574_clk),
    .out(_U574_out)
);
assign _U575_in = _U574_out;
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = _U584_out;
_U576_pt__U577 _U576 (
    .in(_U576_in),
    .out(_U576_out)
);
assign _U578_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U578_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U578 (
    .in(_U578_in),
    .clk(_U578_clk),
    .out(_U578_out)
);
assign _U579_in = _U578_out;
assign _U579_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U579 (
    .in(_U579_in),
    .clk(_U579_clk),
    .out(_U579_out)
);
assign _U580_in = _U579_out;
assign _U580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U580_in),
    .clk(_U580_clk),
    .out(_U580_out)
);
assign _U581_in = _U580_out;
assign _U581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U581_in),
    .clk(_U581_clk),
    .out(_U581_out)
);
assign _U582_in = _U581_out;
assign _U582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U582_in),
    .clk(_U582_clk),
    .out(_U582_out)
);
assign _U583_in = _U582_out;
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = _U583_out;
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign _U585_in = _U593_out;
_U585_pt__U586 _U585 (
    .in(_U585_in),
    .out(_U585_out)
);
assign _U587_in = in1_hw_input_global_wrapper_stencil[7];
assign _U587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U587_in),
    .clk(_U587_clk),
    .out(_U587_out)
);
assign _U588_in = _U587_out;
assign _U588_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(_U588_in),
    .clk(_U588_clk),
    .out(_U588_out)
);
assign _U589_in = _U588_out;
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = _U589_out;
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = _U590_out;
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign _U592_in = _U591_out;
assign _U592_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U592 (
    .in(_U592_in),
    .clk(_U592_clk),
    .out(_U592_out)
);
assign _U593_in = _U592_out;
assign _U593_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U593 (
    .in(_U593_in),
    .clk(_U593_clk),
    .out(_U593_out)
);
assign _U594_in = _U610_out;
_U594_pt__U595 _U594 (
    .in(_U594_in),
    .out(_U594_out)
);
assign _U596_in = 16'(_U506_out * _U508_out);
assign _U596_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U596 (
    .in(_U596_in),
    .clk(_U596_clk),
    .out(_U596_out)
);
assign _U597_in = _U596_out;
assign _U597_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U597 (
    .in(_U597_in),
    .clk(_U597_clk),
    .out(_U597_out)
);
assign _U598_in = _U597_out;
assign _U598_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U598 (
    .in(_U598_in),
    .clk(_U598_clk),
    .out(_U598_out)
);
assign _U599_in = _U598_out;
assign _U599_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U599 (
    .in(_U599_in),
    .clk(_U599_clk),
    .out(_U599_out)
);
assign _U600_in = _U599_out;
assign _U600_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U600 (
    .in(_U600_in),
    .clk(_U600_clk),
    .out(_U600_out)
);
assign _U601_in = _U600_out;
assign _U601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U601_in),
    .clk(_U601_clk),
    .out(_U601_out)
);
assign _U602_in = _U601_out;
assign _U602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U602_in),
    .clk(_U602_clk),
    .out(_U602_out)
);
assign _U603_in = _U602_out;
assign _U603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U603 (
    .in(_U603_in),
    .clk(_U603_clk),
    .out(_U603_out)
);
assign _U604_in = _U603_out;
assign _U604_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U604 (
    .in(_U604_in),
    .clk(_U604_clk),
    .out(_U604_out)
);
assign _U605_in = _U604_out;
assign _U605_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U605 (
    .in(_U605_in),
    .clk(_U605_clk),
    .out(_U605_out)
);
assign _U606_in = _U605_out;
assign _U606_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U606 (
    .in(_U606_in),
    .clk(_U606_clk),
    .out(_U606_out)
);
assign _U607_in = _U606_out;
assign _U607_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U607 (
    .in(_U607_in),
    .clk(_U607_clk),
    .out(_U607_out)
);
assign _U608_in = _U607_out;
assign _U608_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U608 (
    .in(_U608_in),
    .clk(_U608_clk),
    .out(_U608_out)
);
assign _U609_in = _U608_out;
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = _U609_out;
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U408_pt__U409 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_2_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U408_in;
assign _U408_in = 16'h0000;
_U408_pt__U409 _U408 (
    .in(_U408_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U399_pt__U400 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U391_pt__U392 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U383_pt__U384 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U376_pt__U377 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U369_pt__U370 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U363_pt__U364 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U357_pt__U358 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U352_pt__U353 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U347_pt__U348 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U343_pt__U344 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U33_pt__U34 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U339_pt__U340 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U336_pt__U337 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U333_pt__U334 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U331_pt__U332 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U329_pt__U330 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U313_pt__U314 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U310_pt__U311 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U30_pt__U31 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U306_pt__U307 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U303_pt__U304 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U2_pt__U3 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_1_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U2_in;
assign _U2_in = 16'h0000;
_U2_pt__U3 _U2 (
    .in(_U2_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U297_pt__U298 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U294_pt__U295 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U286_pt__U287 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U283_pt__U284 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U27_pt__U28 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U273_pt__U274 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U270_pt__U271 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U258_pt__U259 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U255_pt__U256 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U252_pt__U253 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U238_pt__U239 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U236_pt__U237 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U233_pt__U234 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U216_pt__U217 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U207_pt__U208 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_5_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U207_in;
wire [15:0] _U207_out;
wire [15:0] _U209_in;
wire _U209_clk;
wire [15:0] _U209_out;
wire [15:0] _U210_in;
wire _U210_clk;
wire [15:0] _U210_out;
wire [15:0] _U211_in;
wire _U211_clk;
wire [15:0] _U211_out;
wire [15:0] _U212_in;
wire _U212_clk;
wire [15:0] _U212_out;
wire [15:0] _U213_in;
wire _U213_clk;
wire [15:0] _U213_out;
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire _U215_clk;
wire [15:0] _U215_out;
wire [15:0] _U216_in;
wire [15:0] _U216_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
wire [15:0] _U219_in;
wire _U219_clk;
wire [15:0] _U219_out;
wire [15:0] _U220_in;
wire _U220_clk;
wire [15:0] _U220_out;
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
wire [15:0] _U223_in;
wire _U223_clk;
wire [15:0] _U223_out;
wire [15:0] _U224_in;
wire _U224_clk;
wire [15:0] _U224_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
wire [15:0] _U229_in;
wire _U229_clk;
wire [15:0] _U229_out;
wire [15:0] _U230_in;
wire _U230_clk;
wire [15:0] _U230_out;
wire [15:0] _U231_in;
wire _U231_clk;
wire [15:0] _U231_out;
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
wire [15:0] _U233_in;
wire [15:0] _U233_out;
wire [15:0] _U235_in;
wire _U235_clk;
wire [15:0] _U235_out;
wire [15:0] _U236_in;
wire [15:0] _U238_in;
wire [15:0] _U238_out;
wire [15:0] _U240_in;
wire _U240_clk;
wire [15:0] _U240_out;
wire [15:0] _U241_in;
wire _U241_clk;
wire [15:0] _U241_out;
wire [15:0] _U242_in;
wire _U242_clk;
wire [15:0] _U242_out;
wire [15:0] _U243_in;
wire _U243_clk;
wire [15:0] _U243_out;
wire [15:0] _U244_in;
wire _U244_clk;
wire [15:0] _U244_out;
wire [15:0] _U245_in;
wire _U245_clk;
wire [15:0] _U245_out;
wire [15:0] _U246_in;
wire _U246_clk;
wire [15:0] _U246_out;
wire [15:0] _U247_in;
wire _U247_clk;
wire [15:0] _U247_out;
wire [15:0] _U248_in;
wire _U248_clk;
wire [15:0] _U248_out;
wire [15:0] _U249_in;
wire _U249_clk;
wire [15:0] _U249_out;
wire [15:0] _U250_in;
wire _U250_clk;
wire [15:0] _U250_out;
wire [15:0] _U251_in;
wire _U251_clk;
wire [15:0] _U251_out;
wire [15:0] _U252_in;
wire [15:0] _U252_out;
wire [15:0] _U254_in;
wire _U254_clk;
wire [15:0] _U254_out;
wire [15:0] _U255_in;
wire [15:0] _U255_out;
wire [15:0] _U257_in;
wire _U257_clk;
wire [15:0] _U257_out;
wire [15:0] _U258_in;
wire [15:0] _U258_out;
wire [15:0] _U260_in;
wire _U260_clk;
wire [15:0] _U260_out;
wire [15:0] _U261_in;
wire _U261_clk;
wire [15:0] _U261_out;
wire [15:0] _U262_in;
wire _U262_clk;
wire [15:0] _U262_out;
wire [15:0] _U263_in;
wire _U263_clk;
wire [15:0] _U263_out;
wire [15:0] _U264_in;
wire _U264_clk;
wire [15:0] _U264_out;
wire [15:0] _U265_in;
wire _U265_clk;
wire [15:0] _U265_out;
wire [15:0] _U266_in;
wire _U266_clk;
wire [15:0] _U266_out;
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire _U268_clk;
wire [15:0] _U268_out;
wire [15:0] _U269_in;
wire _U269_clk;
wire [15:0] _U269_out;
wire [15:0] _U270_in;
wire [15:0] _U270_out;
wire [15:0] _U272_in;
wire _U272_clk;
wire [15:0] _U272_out;
wire [15:0] _U273_in;
wire [15:0] _U273_out;
wire [15:0] _U275_in;
wire _U275_clk;
wire [15:0] _U275_out;
wire [15:0] _U276_in;
wire _U276_clk;
wire [15:0] _U276_out;
wire [15:0] _U277_in;
wire _U277_clk;
wire [15:0] _U277_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire _U279_clk;
wire [15:0] _U279_out;
wire [15:0] _U280_in;
wire _U280_clk;
wire [15:0] _U280_out;
wire [15:0] _U281_in;
wire _U281_clk;
wire [15:0] _U281_out;
wire [15:0] _U282_in;
wire _U282_clk;
wire [15:0] _U282_out;
wire [15:0] _U283_in;
wire [15:0] _U283_out;
wire [15:0] _U285_in;
wire _U285_clk;
wire [15:0] _U285_out;
wire [15:0] _U286_in;
wire [15:0] _U286_out;
wire [15:0] _U288_in;
wire _U288_clk;
wire [15:0] _U288_out;
wire [15:0] _U289_in;
wire _U289_clk;
wire [15:0] _U289_out;
wire [15:0] _U290_in;
wire _U290_clk;
wire [15:0] _U290_out;
wire [15:0] _U291_in;
wire _U291_clk;
wire [15:0] _U291_out;
wire [15:0] _U292_in;
wire _U292_clk;
wire [15:0] _U292_out;
wire [15:0] _U293_in;
wire _U293_clk;
wire [15:0] _U293_out;
wire [15:0] _U294_in;
wire [15:0] _U294_out;
wire [15:0] _U296_in;
wire _U296_clk;
wire [15:0] _U296_out;
wire [15:0] _U297_in;
wire [15:0] _U297_out;
wire [15:0] _U299_in;
wire _U299_clk;
wire [15:0] _U299_out;
wire [15:0] _U300_in;
wire _U300_clk;
wire [15:0] _U300_out;
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire [15:0] _U303_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
wire [15:0] _U306_in;
wire [15:0] _U306_out;
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire [15:0] _U310_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
wire [15:0] _U313_in;
wire [15:0] _U313_out;
wire [15:0] _U315_in;
wire _U315_clk;
wire [15:0] _U315_out;
wire [15:0] _U316_in;
wire _U316_clk;
wire [15:0] _U316_out;
wire [15:0] _U317_in;
wire _U317_clk;
wire [15:0] _U317_out;
wire [15:0] _U318_in;
wire _U318_clk;
wire [15:0] _U318_out;
wire [15:0] _U319_in;
wire _U319_clk;
wire [15:0] _U319_out;
wire [15:0] _U320_in;
wire _U320_clk;
wire [15:0] _U320_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire _U322_clk;
wire [15:0] _U322_out;
wire [15:0] _U323_in;
wire _U323_clk;
wire [15:0] _U323_out;
wire [15:0] _U324_in;
wire _U324_clk;
wire [15:0] _U324_out;
wire [15:0] _U325_in;
wire _U325_clk;
wire [15:0] _U325_out;
wire [15:0] _U326_in;
wire _U326_clk;
wire [15:0] _U326_out;
wire [15:0] _U327_in;
wire _U327_clk;
wire [15:0] _U327_out;
wire [15:0] _U328_in;
wire _U328_clk;
wire [15:0] _U328_out;
wire [15:0] _U329_in;
wire [15:0] _U329_out;
wire [15:0] _U331_in;
wire [15:0] _U331_out;
wire [15:0] _U333_in;
wire [15:0] _U333_out;
wire [15:0] _U335_in;
wire _U335_clk;
wire [15:0] _U335_out;
wire [15:0] _U336_in;
wire [15:0] _U336_out;
wire [15:0] _U338_in;
wire _U338_clk;
wire [15:0] _U338_out;
wire [15:0] _U339_in;
wire [15:0] _U339_out;
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire _U342_clk;
wire [15:0] _U342_out;
wire [15:0] _U343_in;
wire [15:0] _U343_out;
wire [15:0] _U345_in;
wire _U345_clk;
wire [15:0] _U345_out;
wire [15:0] _U346_in;
wire _U346_clk;
wire [15:0] _U346_out;
wire [15:0] _U347_in;
wire [15:0] _U347_out;
wire [15:0] _U349_in;
wire _U349_clk;
wire [15:0] _U349_out;
wire [15:0] _U350_in;
wire _U350_clk;
wire [15:0] _U350_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire [15:0] _U352_out;
wire [15:0] _U354_in;
wire _U354_clk;
wire [15:0] _U354_out;
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire _U356_clk;
wire [15:0] _U356_out;
wire [15:0] _U357_in;
wire [15:0] _U357_out;
wire [15:0] _U359_in;
wire _U359_clk;
wire [15:0] _U359_out;
wire [15:0] _U360_in;
wire _U360_clk;
wire [15:0] _U360_out;
wire [15:0] _U361_in;
wire _U361_clk;
wire [15:0] _U361_out;
wire [15:0] _U362_in;
wire _U362_clk;
wire [15:0] _U362_out;
wire [15:0] _U363_in;
wire [15:0] _U363_out;
wire [15:0] _U365_in;
wire _U365_clk;
wire [15:0] _U365_out;
wire [15:0] _U366_in;
wire _U366_clk;
wire [15:0] _U366_out;
wire [15:0] _U367_in;
wire _U367_clk;
wire [15:0] _U367_out;
wire [15:0] _U368_in;
wire _U368_clk;
wire [15:0] _U368_out;
wire [15:0] _U369_in;
wire [15:0] _U369_out;
wire [15:0] _U371_in;
wire _U371_clk;
wire [15:0] _U371_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire _U373_clk;
wire [15:0] _U373_out;
wire [15:0] _U374_in;
wire _U374_clk;
wire [15:0] _U374_out;
wire [15:0] _U375_in;
wire _U375_clk;
wire [15:0] _U375_out;
wire [15:0] _U376_in;
wire [15:0] _U376_out;
wire [15:0] _U378_in;
wire _U378_clk;
wire [15:0] _U378_out;
wire [15:0] _U379_in;
wire _U379_clk;
wire [15:0] _U379_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
wire [15:0] _U381_in;
wire _U381_clk;
wire [15:0] _U381_out;
wire [15:0] _U382_in;
wire _U382_clk;
wire [15:0] _U382_out;
wire [15:0] _U383_in;
wire [15:0] _U383_out;
wire [15:0] _U385_in;
wire _U385_clk;
wire [15:0] _U385_out;
wire [15:0] _U386_in;
wire _U386_clk;
wire [15:0] _U386_out;
wire [15:0] _U387_in;
wire _U387_clk;
wire [15:0] _U387_out;
wire [15:0] _U388_in;
wire _U388_clk;
wire [15:0] _U388_out;
wire [15:0] _U389_in;
wire _U389_clk;
wire [15:0] _U389_out;
wire [15:0] _U390_in;
wire _U390_clk;
wire [15:0] _U390_out;
wire [15:0] _U391_in;
wire [15:0] _U391_out;
wire [15:0] _U393_in;
wire _U393_clk;
wire [15:0] _U393_out;
wire [15:0] _U394_in;
wire _U394_clk;
wire [15:0] _U394_out;
wire [15:0] _U395_in;
wire _U395_clk;
wire [15:0] _U395_out;
wire [15:0] _U396_in;
wire _U396_clk;
wire [15:0] _U396_out;
wire [15:0] _U397_in;
wire _U397_clk;
wire [15:0] _U397_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire [15:0] _U399_out;
wire [15:0] _U401_in;
wire _U401_clk;
wire [15:0] _U401_out;
wire [15:0] _U402_in;
wire _U402_clk;
wire [15:0] _U402_out;
wire [15:0] _U403_in;
wire _U403_clk;
wire [15:0] _U403_out;
wire [15:0] _U404_in;
wire _U404_clk;
wire [15:0] _U404_out;
wire [15:0] _U405_in;
wire _U405_clk;
wire [15:0] _U405_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire _U407_clk;
wire [15:0] _U407_out;
assign _U207_in = _U215_out;
_U207_pt__U208 _U207 (
    .in(_U207_in),
    .out(_U207_out)
);
assign _U209_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U209_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U209 (
    .in(_U209_in),
    .clk(_U209_clk),
    .out(_U209_out)
);
assign _U210_in = _U209_out;
assign _U210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U210 (
    .in(_U210_in),
    .clk(_U210_clk),
    .out(_U210_out)
);
assign _U211_in = _U210_out;
assign _U211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(_U211_in),
    .clk(_U211_clk),
    .out(_U211_out)
);
assign _U212_in = _U211_out;
assign _U212_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U212 (
    .in(_U212_in),
    .clk(_U212_clk),
    .out(_U212_out)
);
assign _U213_in = _U212_out;
assign _U213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(_U213_in),
    .clk(_U213_clk),
    .out(_U213_out)
);
assign _U214_in = _U213_out;
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = _U214_out;
assign _U215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(_U215_in),
    .clk(_U215_clk),
    .out(_U215_out)
);
assign _U216_in = _U232_out;
_U216_pt__U217 _U216 (
    .in(_U216_in),
    .out(_U216_out)
);
assign _U218_in = 16'(_U329_out * _U331_out);
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign _U219_in = _U218_out;
assign _U219_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U219_in),
    .clk(_U219_clk),
    .out(_U219_out)
);
assign _U220_in = _U219_out;
assign _U220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U220_in),
    .clk(_U220_clk),
    .out(_U220_out)
);
assign _U221_in = _U220_out;
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign _U222_in = _U221_out;
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign _U223_in = _U222_out;
assign _U223_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(_U223_in),
    .clk(_U223_clk),
    .out(_U223_out)
);
assign _U224_in = _U223_out;
assign _U224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U224_in),
    .clk(_U224_clk),
    .out(_U224_out)
);
assign _U225_in = _U224_out;
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = _U225_out;
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = _U226_out;
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = _U227_out;
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign _U229_in = _U228_out;
assign _U229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U229_in),
    .clk(_U229_clk),
    .out(_U229_out)
);
assign _U230_in = _U229_out;
assign _U230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U230 (
    .in(_U230_in),
    .clk(_U230_clk),
    .out(_U230_out)
);
assign _U231_in = _U230_out;
assign _U231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U231 (
    .in(_U231_in),
    .clk(_U231_clk),
    .out(_U231_out)
);
assign _U232_in = _U231_out;
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign _U233_in = _U235_out;
_U233_pt__U234 _U233 (
    .in(_U233_in),
    .out(_U233_out)
);
assign _U235_in = 16'(_U313_out + _U255_out);
assign _U235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U235 (
    .in(_U235_in),
    .clk(_U235_clk),
    .out(_U235_out)
);
assign _U236_in = 16'(_U216_out + _U233_out);
_U236_pt__U237 _U236 (
    .in(_U236_in),
    .out(out_conv_stencil)
);
assign _U238_in = _U251_out;
_U238_pt__U239 _U238 (
    .in(_U238_in),
    .out(_U238_out)
);
assign _U240_in = 16'(_U333_out * _U336_out);
assign _U240_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U240 (
    .in(_U240_in),
    .clk(_U240_clk),
    .out(_U240_out)
);
assign _U241_in = _U240_out;
assign _U241_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U241 (
    .in(_U241_in),
    .clk(_U241_clk),
    .out(_U241_out)
);
assign _U242_in = _U241_out;
assign _U242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U242_in),
    .clk(_U242_clk),
    .out(_U242_out)
);
assign _U243_in = _U242_out;
assign _U243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U243_in),
    .clk(_U243_clk),
    .out(_U243_out)
);
assign _U244_in = _U243_out;
assign _U244_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U244 (
    .in(_U244_in),
    .clk(_U244_clk),
    .out(_U244_out)
);
assign _U245_in = _U244_out;
assign _U245_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U245 (
    .in(_U245_in),
    .clk(_U245_clk),
    .out(_U245_out)
);
assign _U246_in = _U245_out;
assign _U246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(_U246_in),
    .clk(_U246_clk),
    .out(_U246_out)
);
assign _U247_in = _U246_out;
assign _U247_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U247 (
    .in(_U247_in),
    .clk(_U247_clk),
    .out(_U247_out)
);
assign _U248_in = _U247_out;
assign _U248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U248 (
    .in(_U248_in),
    .clk(_U248_clk),
    .out(_U248_out)
);
assign _U249_in = _U248_out;
assign _U249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U249 (
    .in(_U249_in),
    .clk(_U249_clk),
    .out(_U249_out)
);
assign _U250_in = _U249_out;
assign _U250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U250 (
    .in(_U250_in),
    .clk(_U250_clk),
    .out(_U250_out)
);
assign _U251_in = _U250_out;
assign _U251_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U251 (
    .in(_U251_in),
    .clk(_U251_clk),
    .out(_U251_out)
);
assign _U252_in = _U254_out;
_U252_pt__U253 _U252 (
    .in(_U252_in),
    .out(_U252_out)
);
assign _U254_in = 16'(_U258_out + _U270_out);
assign _U254_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U254 (
    .in(_U254_in),
    .clk(_U254_clk),
    .out(_U254_out)
);
assign _U255_in = _U257_out;
_U255_pt__U256 _U255 (
    .in(_U255_in),
    .out(_U255_out)
);
assign _U257_in = 16'(_U238_out + _U252_out);
assign _U257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U257 (
    .in(_U257_in),
    .clk(_U257_clk),
    .out(_U257_out)
);
assign _U258_in = _U269_out;
_U258_pt__U259 _U258 (
    .in(_U258_in),
    .out(_U258_out)
);
assign _U260_in = 16'(_U339_out * _U343_out);
assign _U260_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U260_in),
    .clk(_U260_clk),
    .out(_U260_out)
);
assign _U261_in = _U260_out;
assign _U261_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U261 (
    .in(_U261_in),
    .clk(_U261_clk),
    .out(_U261_out)
);
assign _U262_in = _U261_out;
assign _U262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U262 (
    .in(_U262_in),
    .clk(_U262_clk),
    .out(_U262_out)
);
assign _U263_in = _U262_out;
assign _U263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U263 (
    .in(_U263_in),
    .clk(_U263_clk),
    .out(_U263_out)
);
assign _U264_in = _U263_out;
assign _U264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U264_in),
    .clk(_U264_clk),
    .out(_U264_out)
);
assign _U265_in = _U264_out;
assign _U265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U265 (
    .in(_U265_in),
    .clk(_U265_clk),
    .out(_U265_out)
);
assign _U266_in = _U265_out;
assign _U266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U266 (
    .in(_U266_in),
    .clk(_U266_clk),
    .out(_U266_out)
);
assign _U267_in = _U266_out;
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = _U267_out;
assign _U268_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U268 (
    .in(_U268_in),
    .clk(_U268_clk),
    .out(_U268_out)
);
assign _U269_in = _U268_out;
assign _U269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U269 (
    .in(_U269_in),
    .clk(_U269_clk),
    .out(_U269_out)
);
assign _U270_in = _U272_out;
_U270_pt__U271 _U270 (
    .in(_U270_in),
    .out(_U270_out)
);
assign _U272_in = 16'(_U273_out + _U283_out);
assign _U272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U272_in),
    .clk(_U272_clk),
    .out(_U272_out)
);
assign _U273_in = _U282_out;
_U273_pt__U274 _U273 (
    .in(_U273_in),
    .out(_U273_out)
);
assign _U275_in = 16'(_U347_out * _U352_out);
assign _U275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U275 (
    .in(_U275_in),
    .clk(_U275_clk),
    .out(_U275_out)
);
assign _U276_in = _U275_out;
assign _U276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U276 (
    .in(_U276_in),
    .clk(_U276_clk),
    .out(_U276_out)
);
assign _U277_in = _U276_out;
assign _U277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U277 (
    .in(_U277_in),
    .clk(_U277_clk),
    .out(_U277_out)
);
assign _U278_in = _U277_out;
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = _U278_out;
assign _U279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U279_in),
    .clk(_U279_clk),
    .out(_U279_out)
);
assign _U280_in = _U279_out;
assign _U280_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U280 (
    .in(_U280_in),
    .clk(_U280_clk),
    .out(_U280_out)
);
assign _U281_in = _U280_out;
assign _U281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U281_in),
    .clk(_U281_clk),
    .out(_U281_out)
);
assign _U282_in = _U281_out;
assign _U282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U282 (
    .in(_U282_in),
    .clk(_U282_clk),
    .out(_U282_out)
);
assign _U283_in = _U285_out;
_U283_pt__U284 _U283 (
    .in(_U283_in),
    .out(_U283_out)
);
assign _U285_in = 16'(_U286_out + _U294_out);
assign _U285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(_U285_in),
    .clk(_U285_clk),
    .out(_U285_out)
);
assign _U286_in = _U293_out;
_U286_pt__U287 _U286 (
    .in(_U286_in),
    .out(_U286_out)
);
assign _U288_in = 16'(_U357_out * _U363_out);
assign _U288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U288_in),
    .clk(_U288_clk),
    .out(_U288_out)
);
assign _U289_in = _U288_out;
assign _U289_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U289_in),
    .clk(_U289_clk),
    .out(_U289_out)
);
assign _U290_in = _U289_out;
assign _U290_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U290 (
    .in(_U290_in),
    .clk(_U290_clk),
    .out(_U290_out)
);
assign _U291_in = _U290_out;
assign _U291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U291 (
    .in(_U291_in),
    .clk(_U291_clk),
    .out(_U291_out)
);
assign _U292_in = _U291_out;
assign _U292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U292 (
    .in(_U292_in),
    .clk(_U292_clk),
    .out(_U292_out)
);
assign _U293_in = _U292_out;
assign _U293_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U293 (
    .in(_U293_in),
    .clk(_U293_clk),
    .out(_U293_out)
);
assign _U294_in = _U296_out;
_U294_pt__U295 _U294 (
    .in(_U294_in),
    .out(_U294_out)
);
assign _U296_in = 16'(_U297_out + _U303_out);
assign _U296_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U296 (
    .in(_U296_in),
    .clk(_U296_clk),
    .out(_U296_out)
);
assign _U297_in = _U302_out;
_U297_pt__U298 _U297 (
    .in(_U297_in),
    .out(_U297_out)
);
assign _U299_in = 16'(_U369_out * _U376_out);
assign _U299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U299_in),
    .clk(_U299_clk),
    .out(_U299_out)
);
assign _U300_in = _U299_out;
assign _U300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U300 (
    .in(_U300_in),
    .clk(_U300_clk),
    .out(_U300_out)
);
assign _U301_in = _U300_out;
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = _U301_out;
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = _U305_out;
_U303_pt__U304 _U303 (
    .in(_U303_in),
    .out(_U303_out)
);
assign _U305_in = 16'(_U306_out + _U310_out);
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign _U306_in = _U309_out;
_U306_pt__U307 _U306 (
    .in(_U306_in),
    .out(_U306_out)
);
assign _U308_in = 16'(_U383_out * _U391_out);
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = _U308_out;
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = _U312_out;
_U310_pt__U311 _U310 (
    .in(_U310_in),
    .out(_U310_out)
);
assign _U312_in = 16'(_U207_out * _U399_out);
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign _U313_in = _U328_out;
_U313_pt__U314 _U313 (
    .in(_U313_in),
    .out(_U313_out)
);
assign _U315_in = in0_conv_stencil[0];
assign _U315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U315_in),
    .clk(_U315_clk),
    .out(_U315_out)
);
assign _U316_in = _U315_out;
assign _U316_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U316 (
    .in(_U316_in),
    .clk(_U316_clk),
    .out(_U316_out)
);
assign _U317_in = _U316_out;
assign _U317_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U317 (
    .in(_U317_in),
    .clk(_U317_clk),
    .out(_U317_out)
);
assign _U318_in = _U317_out;
assign _U318_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U318 (
    .in(_U318_in),
    .clk(_U318_clk),
    .out(_U318_out)
);
assign _U319_in = _U318_out;
assign _U319_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U319 (
    .in(_U319_in),
    .clk(_U319_clk),
    .out(_U319_out)
);
assign _U320_in = _U319_out;
assign _U320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U320_in),
    .clk(_U320_clk),
    .out(_U320_out)
);
assign _U321_in = _U320_out;
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = _U321_out;
assign _U322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U322 (
    .in(_U322_in),
    .clk(_U322_clk),
    .out(_U322_out)
);
assign _U323_in = _U322_out;
assign _U323_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U323 (
    .in(_U323_in),
    .clk(_U323_clk),
    .out(_U323_out)
);
assign _U324_in = _U323_out;
assign _U324_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U324 (
    .in(_U324_in),
    .clk(_U324_clk),
    .out(_U324_out)
);
assign _U325_in = _U324_out;
assign _U325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U325 (
    .in(_U325_in),
    .clk(_U325_clk),
    .out(_U325_out)
);
assign _U326_in = _U325_out;
assign _U326_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U326 (
    .in(_U326_in),
    .clk(_U326_clk),
    .out(_U326_out)
);
assign _U327_in = _U326_out;
assign _U327_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U327 (
    .in(_U327_in),
    .clk(_U327_clk),
    .out(_U327_out)
);
assign _U328_in = _U327_out;
assign _U328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U328_in),
    .clk(_U328_clk),
    .out(_U328_out)
);
assign _U329_in = in2_hw_kernel_global_wrapper_stencil[0];
_U329_pt__U330 _U329 (
    .in(_U329_in),
    .out(_U329_out)
);
assign _U331_in = in1_hw_input_global_wrapper_stencil[0];
_U331_pt__U332 _U331 (
    .in(_U331_in),
    .out(_U331_out)
);
assign _U333_in = _U335_out;
_U333_pt__U334 _U333 (
    .in(_U333_in),
    .out(_U333_out)
);
assign _U335_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U335 (
    .in(_U335_in),
    .clk(_U335_clk),
    .out(_U335_out)
);
assign _U336_in = _U338_out;
_U336_pt__U337 _U336 (
    .in(_U336_in),
    .out(_U336_out)
);
assign _U338_in = in1_hw_input_global_wrapper_stencil[1];
assign _U338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U338_in),
    .clk(_U338_clk),
    .out(_U338_out)
);
assign _U339_in = _U342_out;
_U339_pt__U340 _U339 (
    .in(_U339_in),
    .out(_U339_out)
);
assign _U341_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = _U341_out;
assign _U342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U342_in),
    .clk(_U342_clk),
    .out(_U342_out)
);
assign _U343_in = _U346_out;
_U343_pt__U344 _U343 (
    .in(_U343_in),
    .out(_U343_out)
);
assign _U345_in = in1_hw_input_global_wrapper_stencil[2];
assign _U345_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(_U345_in),
    .clk(_U345_clk),
    .out(_U345_out)
);
assign _U346_in = _U345_out;
assign _U346_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U346 (
    .in(_U346_in),
    .clk(_U346_clk),
    .out(_U346_out)
);
assign _U347_in = _U351_out;
_U347_pt__U348 _U347 (
    .in(_U347_in),
    .out(_U347_out)
);
assign _U349_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U349_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U349 (
    .in(_U349_in),
    .clk(_U349_clk),
    .out(_U349_out)
);
assign _U350_in = _U349_out;
assign _U350_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U350_in),
    .clk(_U350_clk),
    .out(_U350_out)
);
assign _U351_in = _U350_out;
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = _U356_out;
_U352_pt__U353 _U352 (
    .in(_U352_in),
    .out(_U352_out)
);
assign _U354_in = in1_hw_input_global_wrapper_stencil[3];
assign _U354_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U354 (
    .in(_U354_in),
    .clk(_U354_clk),
    .out(_U354_out)
);
assign _U355_in = _U354_out;
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = _U355_out;
assign _U356_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U356 (
    .in(_U356_in),
    .clk(_U356_clk),
    .out(_U356_out)
);
assign _U357_in = _U362_out;
_U357_pt__U358 _U357 (
    .in(_U357_in),
    .out(_U357_out)
);
assign _U359_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U359 (
    .in(_U359_in),
    .clk(_U359_clk),
    .out(_U359_out)
);
assign _U360_in = _U359_out;
assign _U360_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U360 (
    .in(_U360_in),
    .clk(_U360_clk),
    .out(_U360_out)
);
assign _U361_in = _U360_out;
assign _U361_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U361 (
    .in(_U361_in),
    .clk(_U361_clk),
    .out(_U361_out)
);
assign _U362_in = _U361_out;
assign _U362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U362 (
    .in(_U362_in),
    .clk(_U362_clk),
    .out(_U362_out)
);
assign _U363_in = _U368_out;
_U363_pt__U364 _U363 (
    .in(_U363_in),
    .out(_U363_out)
);
assign _U365_in = in1_hw_input_global_wrapper_stencil[4];
assign _U365_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U365 (
    .in(_U365_in),
    .clk(_U365_clk),
    .out(_U365_out)
);
assign _U366_in = _U365_out;
assign _U366_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U366 (
    .in(_U366_in),
    .clk(_U366_clk),
    .out(_U366_out)
);
assign _U367_in = _U366_out;
assign _U367_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U367 (
    .in(_U367_in),
    .clk(_U367_clk),
    .out(_U367_out)
);
assign _U368_in = _U367_out;
assign _U368_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U368 (
    .in(_U368_in),
    .clk(_U368_clk),
    .out(_U368_out)
);
assign _U369_in = _U375_out;
_U369_pt__U370 _U369 (
    .in(_U369_in),
    .out(_U369_out)
);
assign _U371_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U371_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(_U371_in),
    .clk(_U371_clk),
    .out(_U371_out)
);
assign _U372_in = _U371_out;
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = _U372_out;
assign _U373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U373 (
    .in(_U373_in),
    .clk(_U373_clk),
    .out(_U373_out)
);
assign _U374_in = _U373_out;
assign _U374_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U374 (
    .in(_U374_in),
    .clk(_U374_clk),
    .out(_U374_out)
);
assign _U375_in = _U374_out;
assign _U375_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U375 (
    .in(_U375_in),
    .clk(_U375_clk),
    .out(_U375_out)
);
assign _U376_in = _U382_out;
_U376_pt__U377 _U376 (
    .in(_U376_in),
    .out(_U376_out)
);
assign _U378_in = in1_hw_input_global_wrapper_stencil[5];
assign _U378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U378_in),
    .clk(_U378_clk),
    .out(_U378_out)
);
assign _U379_in = _U378_out;
assign _U379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U379_in),
    .clk(_U379_clk),
    .out(_U379_out)
);
assign _U380_in = _U379_out;
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign _U381_in = _U380_out;
assign _U381_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U381 (
    .in(_U381_in),
    .clk(_U381_clk),
    .out(_U381_out)
);
assign _U382_in = _U381_out;
assign _U382_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U382 (
    .in(_U382_in),
    .clk(_U382_clk),
    .out(_U382_out)
);
assign _U383_in = _U390_out;
_U383_pt__U384 _U383 (
    .in(_U383_in),
    .out(_U383_out)
);
assign _U385_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U385_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U385 (
    .in(_U385_in),
    .clk(_U385_clk),
    .out(_U385_out)
);
assign _U386_in = _U385_out;
assign _U386_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U386 (
    .in(_U386_in),
    .clk(_U386_clk),
    .out(_U386_out)
);
assign _U387_in = _U386_out;
assign _U387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U387 (
    .in(_U387_in),
    .clk(_U387_clk),
    .out(_U387_out)
);
assign _U388_in = _U387_out;
assign _U388_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U388 (
    .in(_U388_in),
    .clk(_U388_clk),
    .out(_U388_out)
);
assign _U389_in = _U388_out;
assign _U389_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U389 (
    .in(_U389_in),
    .clk(_U389_clk),
    .out(_U389_out)
);
assign _U390_in = _U389_out;
assign _U390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(_U390_in),
    .clk(_U390_clk),
    .out(_U390_out)
);
assign _U391_in = _U398_out;
_U391_pt__U392 _U391 (
    .in(_U391_in),
    .out(_U391_out)
);
assign _U393_in = in1_hw_input_global_wrapper_stencil[6];
assign _U393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U393 (
    .in(_U393_in),
    .clk(_U393_clk),
    .out(_U393_out)
);
assign _U394_in = _U393_out;
assign _U394_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U394 (
    .in(_U394_in),
    .clk(_U394_clk),
    .out(_U394_out)
);
assign _U395_in = _U394_out;
assign _U395_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U395 (
    .in(_U395_in),
    .clk(_U395_clk),
    .out(_U395_out)
);
assign _U396_in = _U395_out;
assign _U396_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U396 (
    .in(_U396_in),
    .clk(_U396_clk),
    .out(_U396_out)
);
assign _U397_in = _U396_out;
assign _U397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U397_in),
    .clk(_U397_clk),
    .out(_U397_out)
);
assign _U398_in = _U397_out;
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = _U407_out;
_U399_pt__U400 _U399 (
    .in(_U399_in),
    .out(_U399_out)
);
assign _U401_in = in1_hw_input_global_wrapper_stencil[7];
assign _U401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U401_in),
    .clk(_U401_clk),
    .out(_U401_out)
);
assign _U402_in = _U401_out;
assign _U402_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U402 (
    .in(_U402_in),
    .clk(_U402_clk),
    .out(_U402_out)
);
assign _U403_in = _U402_out;
assign _U403_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U403 (
    .in(_U403_in),
    .clk(_U403_clk),
    .out(_U403_out)
);
assign _U404_in = _U403_out;
assign _U404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U404 (
    .in(_U404_in),
    .clk(_U404_clk),
    .out(_U404_out)
);
assign _U405_in = _U404_out;
assign _U405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(_U405_in),
    .clk(_U405_clk),
    .out(_U405_out)
);
assign _U406_in = _U405_out;
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = _U406_out;
assign _U407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U407 (
    .in(_U407_in),
    .clk(_U407_clk),
    .out(_U407_out)
);
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U205_pt__U206 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U205_in;
assign _U205_in = 16'h0000;
_U205_pt__U206 _U205 (
    .in(_U205_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U189_pt__U190 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U173_pt__U174 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U165_pt__U166 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U157_pt__U158 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U150_pt__U151 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U143_pt__U144 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U13_pt__U14 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U137_pt__U138 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U131_pt__U132 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U126_pt__U127 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U121_pt__U122 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U11_pt__U12 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U117_pt__U118 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U113_pt__U114 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U110_pt__U111 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U107_pt__U108 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U105_pt__U106 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U103_pt__U104 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_4_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U10_in;
wire _U10_clk;
wire [15:0] _U10_out;
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U102_in;
wire _U102_clk;
wire [15:0] _U102_out;
wire [15:0] _U103_in;
wire [15:0] _U103_out;
wire [15:0] _U105_in;
wire [15:0] _U105_out;
wire [15:0] _U107_in;
wire [15:0] _U107_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
wire [15:0] _U11_in;
wire [15:0] _U110_in;
wire [15:0] _U110_out;
wire [15:0] _U112_in;
wire _U112_clk;
wire [15:0] _U112_out;
wire [15:0] _U113_in;
wire [15:0] _U113_out;
wire [15:0] _U115_in;
wire _U115_clk;
wire [15:0] _U115_out;
wire [15:0] _U116_in;
wire _U116_clk;
wire [15:0] _U116_out;
wire [15:0] _U117_in;
wire [15:0] _U117_out;
wire [15:0] _U119_in;
wire _U119_clk;
wire [15:0] _U119_out;
wire [15:0] _U120_in;
wire _U120_clk;
wire [15:0] _U120_out;
wire [15:0] _U121_in;
wire [15:0] _U121_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
wire [15:0] _U125_in;
wire _U125_clk;
wire [15:0] _U125_out;
wire [15:0] _U126_in;
wire [15:0] _U126_out;
wire [15:0] _U128_in;
wire _U128_clk;
wire [15:0] _U128_out;
wire [15:0] _U129_in;
wire _U129_clk;
wire [15:0] _U129_out;
wire [15:0] _U13_in;
wire [15:0] _U13_out;
wire [15:0] _U130_in;
wire _U130_clk;
wire [15:0] _U130_out;
wire [15:0] _U131_in;
wire [15:0] _U131_out;
wire [15:0] _U133_in;
wire _U133_clk;
wire [15:0] _U133_out;
wire [15:0] _U134_in;
wire _U134_clk;
wire [15:0] _U134_out;
wire [15:0] _U135_in;
wire _U135_clk;
wire [15:0] _U135_out;
wire [15:0] _U136_in;
wire _U136_clk;
wire [15:0] _U136_out;
wire [15:0] _U137_in;
wire [15:0] _U137_out;
wire [15:0] _U139_in;
wire _U139_clk;
wire [15:0] _U139_out;
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire _U141_clk;
wire [15:0] _U141_out;
wire [15:0] _U142_in;
wire _U142_clk;
wire [15:0] _U142_out;
wire [15:0] _U143_in;
wire [15:0] _U143_out;
wire [15:0] _U145_in;
wire _U145_clk;
wire [15:0] _U145_out;
wire [15:0] _U146_in;
wire _U146_clk;
wire [15:0] _U146_out;
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire _U148_clk;
wire [15:0] _U148_out;
wire [15:0] _U149_in;
wire _U149_clk;
wire [15:0] _U149_out;
wire [15:0] _U15_in;
wire _U15_clk;
wire [15:0] _U15_out;
wire [15:0] _U150_in;
wire [15:0] _U150_out;
wire [15:0] _U152_in;
wire _U152_clk;
wire [15:0] _U152_out;
wire [15:0] _U153_in;
wire _U153_clk;
wire [15:0] _U153_out;
wire [15:0] _U154_in;
wire _U154_clk;
wire [15:0] _U154_out;
wire [15:0] _U155_in;
wire _U155_clk;
wire [15:0] _U155_out;
wire [15:0] _U156_in;
wire _U156_clk;
wire [15:0] _U156_out;
wire [15:0] _U157_in;
wire [15:0] _U157_out;
wire [15:0] _U159_in;
wire _U159_clk;
wire [15:0] _U159_out;
wire [15:0] _U16_in;
wire _U16_clk;
wire [15:0] _U16_out;
wire [15:0] _U160_in;
wire _U160_clk;
wire [15:0] _U160_out;
wire [15:0] _U161_in;
wire _U161_clk;
wire [15:0] _U161_out;
wire [15:0] _U162_in;
wire _U162_clk;
wire [15:0] _U162_out;
wire [15:0] _U163_in;
wire _U163_clk;
wire [15:0] _U163_out;
wire [15:0] _U164_in;
wire _U164_clk;
wire [15:0] _U164_out;
wire [15:0] _U165_in;
wire [15:0] _U165_out;
wire [15:0] _U167_in;
wire _U167_clk;
wire [15:0] _U167_out;
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
wire [15:0] _U169_in;
wire _U169_clk;
wire [15:0] _U169_out;
wire [15:0] _U17_in;
wire _U17_clk;
wire [15:0] _U17_out;
wire [15:0] _U170_in;
wire _U170_clk;
wire [15:0] _U170_out;
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire _U172_clk;
wire [15:0] _U172_out;
wire [15:0] _U173_in;
wire [15:0] _U173_out;
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
wire [15:0] _U176_in;
wire _U176_clk;
wire [15:0] _U176_out;
wire [15:0] _U177_in;
wire _U177_clk;
wire [15:0] _U177_out;
wire [15:0] _U178_in;
wire _U178_clk;
wire [15:0] _U178_out;
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
wire [15:0] _U18_in;
wire _U18_clk;
wire [15:0] _U18_out;
wire [15:0] _U180_in;
wire _U180_clk;
wire [15:0] _U180_out;
wire [15:0] _U181_in;
wire _U181_clk;
wire [15:0] _U181_out;
wire [15:0] _U182_in;
wire _U182_clk;
wire [15:0] _U182_out;
wire [15:0] _U183_in;
wire _U183_clk;
wire [15:0] _U183_out;
wire [15:0] _U184_in;
wire _U184_clk;
wire [15:0] _U184_out;
wire [15:0] _U185_in;
wire _U185_clk;
wire [15:0] _U185_out;
wire [15:0] _U186_in;
wire _U186_clk;
wire [15:0] _U186_out;
wire [15:0] _U187_in;
wire _U187_clk;
wire [15:0] _U187_out;
wire [15:0] _U188_in;
wire _U188_clk;
wire [15:0] _U188_out;
wire [15:0] _U189_in;
wire [15:0] _U189_out;
wire [15:0] _U19_in;
wire _U19_clk;
wire [15:0] _U19_out;
wire [15:0] _U191_in;
wire _U191_clk;
wire [15:0] _U191_out;
wire [15:0] _U192_in;
wire _U192_clk;
wire [15:0] _U192_out;
wire [15:0] _U193_in;
wire _U193_clk;
wire [15:0] _U193_out;
wire [15:0] _U194_in;
wire _U194_clk;
wire [15:0] _U194_out;
wire [15:0] _U195_in;
wire _U195_clk;
wire [15:0] _U195_out;
wire [15:0] _U196_in;
wire _U196_clk;
wire [15:0] _U196_out;
wire [15:0] _U197_in;
wire _U197_clk;
wire [15:0] _U197_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire _U199_clk;
wire [15:0] _U199_out;
wire [15:0] _U20_in;
wire _U20_clk;
wire [15:0] _U20_out;
wire [15:0] _U200_in;
wire _U200_clk;
wire [15:0] _U200_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
wire [15:0] _U202_in;
wire _U202_clk;
wire [15:0] _U202_out;
wire [15:0] _U203_in;
wire _U203_clk;
wire [15:0] _U203_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U21_in;
wire _U21_clk;
wire [15:0] _U21_out;
wire [15:0] _U22_in;
wire _U22_clk;
wire [15:0] _U22_out;
wire [15:0] _U23_in;
wire _U23_clk;
wire [15:0] _U23_out;
wire [15:0] _U24_in;
wire _U24_clk;
wire [15:0] _U24_out;
wire [15:0] _U25_in;
wire _U25_clk;
wire [15:0] _U25_out;
wire [15:0] _U26_in;
wire _U26_clk;
wire [15:0] _U26_out;
wire [15:0] _U27_in;
wire [15:0] _U27_out;
wire [15:0] _U29_in;
wire _U29_clk;
wire [15:0] _U29_out;
wire [15:0] _U30_in;
wire [15:0] _U30_out;
wire [15:0] _U32_in;
wire _U32_clk;
wire [15:0] _U32_out;
wire [15:0] _U33_in;
wire [15:0] _U33_out;
wire [15:0] _U35_in;
wire _U35_clk;
wire [15:0] _U35_out;
wire [15:0] _U36_in;
wire _U36_clk;
wire [15:0] _U36_out;
wire [15:0] _U37_in;
wire _U37_clk;
wire [15:0] _U37_out;
wire [15:0] _U38_in;
wire _U38_clk;
wire [15:0] _U38_out;
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
wire [15:0] _U4_in;
wire [15:0] _U4_out;
wire [15:0] _U40_in;
wire _U40_clk;
wire [15:0] _U40_out;
wire [15:0] _U41_in;
wire _U41_clk;
wire [15:0] _U41_out;
wire [15:0] _U42_in;
wire _U42_clk;
wire [15:0] _U42_out;
wire [15:0] _U43_in;
wire _U43_clk;
wire [15:0] _U43_out;
wire [15:0] _U44_in;
wire _U44_clk;
wire [15:0] _U44_out;
wire [15:0] _U45_in;
wire [15:0] _U45_out;
wire [15:0] _U47_in;
wire _U47_clk;
wire [15:0] _U47_out;
wire [15:0] _U48_in;
wire [15:0] _U48_out;
wire [15:0] _U50_in;
wire _U50_clk;
wire [15:0] _U50_out;
wire [15:0] _U51_in;
wire _U51_clk;
wire [15:0] _U51_out;
wire [15:0] _U52_in;
wire _U52_clk;
wire [15:0] _U52_out;
wire [15:0] _U53_in;
wire _U53_clk;
wire [15:0] _U53_out;
wire [15:0] _U54_in;
wire _U54_clk;
wire [15:0] _U54_out;
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
wire [15:0] _U56_in;
wire _U56_clk;
wire [15:0] _U56_out;
wire [15:0] _U57_in;
wire _U57_clk;
wire [15:0] _U57_out;
wire [15:0] _U58_in;
wire [15:0] _U58_out;
wire [15:0] _U6_in;
wire _U6_clk;
wire [15:0] _U6_out;
wire [15:0] _U60_in;
wire _U60_clk;
wire [15:0] _U60_out;
wire [15:0] _U61_in;
wire [15:0] _U61_out;
wire [15:0] _U63_in;
wire _U63_clk;
wire [15:0] _U63_out;
wire [15:0] _U64_in;
wire _U64_clk;
wire [15:0] _U64_out;
wire [15:0] _U65_in;
wire _U65_clk;
wire [15:0] _U65_out;
wire [15:0] _U66_in;
wire _U66_clk;
wire [15:0] _U66_out;
wire [15:0] _U67_in;
wire _U67_clk;
wire [15:0] _U67_out;
wire [15:0] _U68_in;
wire _U68_clk;
wire [15:0] _U68_out;
wire [15:0] _U69_in;
wire [15:0] _U69_out;
wire [15:0] _U7_in;
wire [15:0] _U7_out;
wire [15:0] _U71_in;
wire _U71_clk;
wire [15:0] _U71_out;
wire [15:0] _U72_in;
wire [15:0] _U72_out;
wire [15:0] _U74_in;
wire _U74_clk;
wire [15:0] _U74_out;
wire [15:0] _U75_in;
wire _U75_clk;
wire [15:0] _U75_out;
wire [15:0] _U76_in;
wire _U76_clk;
wire [15:0] _U76_out;
wire [15:0] _U77_in;
wire _U77_clk;
wire [15:0] _U77_out;
wire [15:0] _U78_in;
wire [15:0] _U78_out;
wire [15:0] _U80_in;
wire _U80_clk;
wire [15:0] _U80_out;
wire [15:0] _U81_in;
wire [15:0] _U81_out;
wire [15:0] _U83_in;
wire _U83_clk;
wire [15:0] _U83_out;
wire [15:0] _U84_in;
wire _U84_clk;
wire [15:0] _U84_out;
wire [15:0] _U85_in;
wire [15:0] _U85_out;
wire [15:0] _U87_in;
wire _U87_clk;
wire [15:0] _U87_out;
wire [15:0] _U88_in;
wire [15:0] _U88_out;
wire [15:0] _U9_in;
wire _U9_clk;
wire [15:0] _U9_out;
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
wire [15:0] _U93_in;
wire _U93_clk;
wire [15:0] _U93_out;
wire [15:0] _U94_in;
wire _U94_clk;
wire [15:0] _U94_out;
wire [15:0] _U95_in;
wire _U95_clk;
wire [15:0] _U95_out;
wire [15:0] _U96_in;
wire _U96_clk;
wire [15:0] _U96_out;
wire [15:0] _U97_in;
wire _U97_clk;
wire [15:0] _U97_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U10_in = _U9_out;
assign _U10_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U10 (
    .in(_U10_in),
    .clk(_U10_clk),
    .out(_U10_out)
);
assign _U100_in = _U99_out;
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = _U100_out;
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U102_in = _U101_out;
assign _U102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U102_in),
    .clk(_U102_clk),
    .out(_U102_out)
);
assign _U103_in = in2_hw_kernel_global_wrapper_stencil[0];
_U103_pt__U104 _U103 (
    .in(_U103_in),
    .out(_U103_out)
);
assign _U105_in = in1_hw_input_global_wrapper_stencil[0];
_U105_pt__U106 _U105 (
    .in(_U105_in),
    .out(_U105_out)
);
assign _U107_in = _U109_out;
_U107_pt__U108 _U107 (
    .in(_U107_in),
    .out(_U107_out)
);
assign _U109_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign _U11_in = 16'(_U4_out + _U7_out);
_U11_pt__U12 _U11 (
    .in(_U11_in),
    .out(out_conv_stencil)
);
assign _U110_in = _U112_out;
_U110_pt__U111 _U110 (
    .in(_U110_in),
    .out(_U110_out)
);
assign _U112_in = in1_hw_input_global_wrapper_stencil[1];
assign _U112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U112_in),
    .clk(_U112_clk),
    .out(_U112_out)
);
assign _U113_in = _U116_out;
_U113_pt__U114 _U113 (
    .in(_U113_in),
    .out(_U113_out)
);
assign _U115_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U115_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U115 (
    .in(_U115_in),
    .clk(_U115_clk),
    .out(_U115_out)
);
assign _U116_in = _U115_out;
assign _U116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U116_in),
    .clk(_U116_clk),
    .out(_U116_out)
);
assign _U117_in = _U120_out;
_U117_pt__U118 _U117 (
    .in(_U117_in),
    .out(_U117_out)
);
assign _U119_in = in1_hw_input_global_wrapper_stencil[2];
assign _U119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U119 (
    .in(_U119_in),
    .clk(_U119_clk),
    .out(_U119_out)
);
assign _U120_in = _U119_out;
assign _U120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(_U120_in),
    .clk(_U120_clk),
    .out(_U120_out)
);
assign _U121_in = _U125_out;
_U121_pt__U122 _U121 (
    .in(_U121_in),
    .out(_U121_out)
);
assign _U123_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = _U123_out;
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign _U125_in = _U124_out;
assign _U125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U125 (
    .in(_U125_in),
    .clk(_U125_clk),
    .out(_U125_out)
);
assign _U126_in = _U130_out;
_U126_pt__U127 _U126 (
    .in(_U126_in),
    .out(_U126_out)
);
assign _U128_in = in1_hw_input_global_wrapper_stencil[3];
assign _U128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U128_in),
    .clk(_U128_clk),
    .out(_U128_out)
);
assign _U129_in = _U128_out;
assign _U129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U129_in),
    .clk(_U129_clk),
    .out(_U129_out)
);
assign _U13_in = _U26_out;
_U13_pt__U14 _U13 (
    .in(_U13_in),
    .out(_U13_out)
);
assign _U130_in = _U129_out;
assign _U130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U130_in),
    .clk(_U130_clk),
    .out(_U130_out)
);
assign _U131_in = _U136_out;
_U131_pt__U132 _U131 (
    .in(_U131_in),
    .out(_U131_out)
);
assign _U133_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U133_in),
    .clk(_U133_clk),
    .out(_U133_out)
);
assign _U134_in = _U133_out;
assign _U134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U134_in),
    .clk(_U134_clk),
    .out(_U134_out)
);
assign _U135_in = _U134_out;
assign _U135_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U135 (
    .in(_U135_in),
    .clk(_U135_clk),
    .out(_U135_out)
);
assign _U136_in = _U135_out;
assign _U136_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U136 (
    .in(_U136_in),
    .clk(_U136_clk),
    .out(_U136_out)
);
assign _U137_in = _U142_out;
_U137_pt__U138 _U137 (
    .in(_U137_in),
    .out(_U137_out)
);
assign _U139_in = in1_hw_input_global_wrapper_stencil[4];
assign _U139_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U139 (
    .in(_U139_in),
    .clk(_U139_clk),
    .out(_U139_out)
);
assign _U140_in = _U139_out;
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = _U140_out;
assign _U141_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U141 (
    .in(_U141_in),
    .clk(_U141_clk),
    .out(_U141_out)
);
assign _U142_in = _U141_out;
assign _U142_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U142 (
    .in(_U142_in),
    .clk(_U142_clk),
    .out(_U142_out)
);
assign _U143_in = _U149_out;
_U143_pt__U144 _U143 (
    .in(_U143_in),
    .out(_U143_out)
);
assign _U145_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U145_in),
    .clk(_U145_clk),
    .out(_U145_out)
);
assign _U146_in = _U145_out;
assign _U146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U146_in),
    .clk(_U146_clk),
    .out(_U146_out)
);
assign _U147_in = _U146_out;
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = _U147_out;
assign _U148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U148_in),
    .clk(_U148_clk),
    .out(_U148_out)
);
assign _U149_in = _U148_out;
assign _U149_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U149 (
    .in(_U149_in),
    .clk(_U149_clk),
    .out(_U149_out)
);
assign _U15_in = 16'(_U103_out * _U105_out);
assign _U15_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U15 (
    .in(_U15_in),
    .clk(_U15_clk),
    .out(_U15_out)
);
assign _U150_in = _U156_out;
_U150_pt__U151 _U150 (
    .in(_U150_in),
    .out(_U150_out)
);
assign _U152_in = in1_hw_input_global_wrapper_stencil[5];
assign _U152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U152 (
    .in(_U152_in),
    .clk(_U152_clk),
    .out(_U152_out)
);
assign _U153_in = _U152_out;
assign _U153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U153 (
    .in(_U153_in),
    .clk(_U153_clk),
    .out(_U153_out)
);
assign _U154_in = _U153_out;
assign _U154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(_U154_in),
    .clk(_U154_clk),
    .out(_U154_out)
);
assign _U155_in = _U154_out;
assign _U155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U155_in),
    .clk(_U155_clk),
    .out(_U155_out)
);
assign _U156_in = _U155_out;
assign _U156_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U156 (
    .in(_U156_in),
    .clk(_U156_clk),
    .out(_U156_out)
);
assign _U157_in = _U164_out;
_U157_pt__U158 _U157 (
    .in(_U157_in),
    .out(_U157_out)
);
assign _U159_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U159_in),
    .clk(_U159_clk),
    .out(_U159_out)
);
assign _U16_in = _U15_out;
assign _U16_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U16 (
    .in(_U16_in),
    .clk(_U16_clk),
    .out(_U16_out)
);
assign _U160_in = _U159_out;
assign _U160_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U160 (
    .in(_U160_in),
    .clk(_U160_clk),
    .out(_U160_out)
);
assign _U161_in = _U160_out;
assign _U161_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U161 (
    .in(_U161_in),
    .clk(_U161_clk),
    .out(_U161_out)
);
assign _U162_in = _U161_out;
assign _U162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(_U162_in),
    .clk(_U162_clk),
    .out(_U162_out)
);
assign _U163_in = _U162_out;
assign _U163_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(_U163_in),
    .clk(_U163_clk),
    .out(_U163_out)
);
assign _U164_in = _U163_out;
assign _U164_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(_U164_in),
    .clk(_U164_clk),
    .out(_U164_out)
);
assign _U165_in = _U172_out;
_U165_pt__U166 _U165 (
    .in(_U165_in),
    .out(_U165_out)
);
assign _U167_in = in1_hw_input_global_wrapper_stencil[6];
assign _U167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U167_in),
    .clk(_U167_clk),
    .out(_U167_out)
);
assign _U168_in = _U167_out;
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign _U169_in = _U168_out;
assign _U169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U169 (
    .in(_U169_in),
    .clk(_U169_clk),
    .out(_U169_out)
);
assign _U17_in = _U16_out;
assign _U17_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U17 (
    .in(_U17_in),
    .clk(_U17_clk),
    .out(_U17_out)
);
assign _U170_in = _U169_out;
assign _U170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U170 (
    .in(_U170_in),
    .clk(_U170_clk),
    .out(_U170_out)
);
assign _U171_in = _U170_out;
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = _U171_out;
assign _U172_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(_U172_in),
    .clk(_U172_clk),
    .out(_U172_out)
);
assign _U173_in = _U188_out;
_U173_pt__U174 _U173 (
    .in(_U173_in),
    .out(_U173_out)
);
assign _U175_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign _U176_in = _U175_out;
assign _U176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U176 (
    .in(_U176_in),
    .clk(_U176_clk),
    .out(_U176_out)
);
assign _U177_in = _U176_out;
assign _U177_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U177 (
    .in(_U177_in),
    .clk(_U177_clk),
    .out(_U177_out)
);
assign _U178_in = _U177_out;
assign _U178_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U178 (
    .in(_U178_in),
    .clk(_U178_clk),
    .out(_U178_out)
);
assign _U179_in = _U178_out;
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign _U18_in = _U17_out;
assign _U18_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U18 (
    .in(_U18_in),
    .clk(_U18_clk),
    .out(_U18_out)
);
assign _U180_in = _U179_out;
assign _U180_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U180 (
    .in(_U180_in),
    .clk(_U180_clk),
    .out(_U180_out)
);
assign _U181_in = _U180_out;
assign _U181_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U181 (
    .in(_U181_in),
    .clk(_U181_clk),
    .out(_U181_out)
);
assign _U182_in = _U181_out;
assign _U182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U182_in),
    .clk(_U182_clk),
    .out(_U182_out)
);
assign _U183_in = _U182_out;
assign _U183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U183_in),
    .clk(_U183_clk),
    .out(_U183_out)
);
assign _U184_in = _U183_out;
assign _U184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U184_in),
    .clk(_U184_clk),
    .out(_U184_out)
);
assign _U185_in = _U184_out;
assign _U185_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U185 (
    .in(_U185_in),
    .clk(_U185_clk),
    .out(_U185_out)
);
assign _U186_in = _U185_out;
assign _U186_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U186 (
    .in(_U186_in),
    .clk(_U186_clk),
    .out(_U186_out)
);
assign _U187_in = _U186_out;
assign _U187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U187 (
    .in(_U187_in),
    .clk(_U187_clk),
    .out(_U187_out)
);
assign _U188_in = _U187_out;
assign _U188_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U188 (
    .in(_U188_in),
    .clk(_U188_clk),
    .out(_U188_out)
);
assign _U189_in = _U204_out;
_U189_pt__U190 _U189 (
    .in(_U189_in),
    .out(_U189_out)
);
assign _U19_in = _U18_out;
assign _U19_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U19 (
    .in(_U19_in),
    .clk(_U19_clk),
    .out(_U19_out)
);
assign _U191_in = in1_hw_input_global_wrapper_stencil[7];
assign _U191_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U191_in),
    .clk(_U191_clk),
    .out(_U191_out)
);
assign _U192_in = _U191_out;
assign _U192_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U192_in),
    .clk(_U192_clk),
    .out(_U192_out)
);
assign _U193_in = _U192_out;
assign _U193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U193_in),
    .clk(_U193_clk),
    .out(_U193_out)
);
assign _U194_in = _U193_out;
assign _U194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U194 (
    .in(_U194_in),
    .clk(_U194_clk),
    .out(_U194_out)
);
assign _U195_in = _U194_out;
assign _U195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U195 (
    .in(_U195_in),
    .clk(_U195_clk),
    .out(_U195_out)
);
assign _U196_in = _U195_out;
assign _U196_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U196 (
    .in(_U196_in),
    .clk(_U196_clk),
    .out(_U196_out)
);
assign _U197_in = _U196_out;
assign _U197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U197 (
    .in(_U197_in),
    .clk(_U197_clk),
    .out(_U197_out)
);
assign _U198_in = _U197_out;
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = _U198_out;
assign _U199_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U199 (
    .in(_U199_in),
    .clk(_U199_clk),
    .out(_U199_out)
);
assign _U20_in = _U19_out;
assign _U20_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U20 (
    .in(_U20_in),
    .clk(_U20_clk),
    .out(_U20_out)
);
assign _U200_in = _U199_out;
assign _U200_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U200 (
    .in(_U200_in),
    .clk(_U200_clk),
    .out(_U200_out)
);
assign _U201_in = _U200_out;
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign _U202_in = _U201_out;
assign _U202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U202 (
    .in(_U202_in),
    .clk(_U202_clk),
    .out(_U202_out)
);
assign _U203_in = _U202_out;
assign _U203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U203 (
    .in(_U203_in),
    .clk(_U203_clk),
    .out(_U203_out)
);
assign _U204_in = _U203_out;
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U21_in = _U20_out;
assign _U21_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U21 (
    .in(_U21_in),
    .clk(_U21_clk),
    .out(_U21_out)
);
assign _U22_in = _U21_out;
assign _U22_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U22 (
    .in(_U22_in),
    .clk(_U22_clk),
    .out(_U22_out)
);
assign _U23_in = _U22_out;
assign _U23_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U23 (
    .in(_U23_in),
    .clk(_U23_clk),
    .out(_U23_out)
);
assign _U24_in = _U23_out;
assign _U24_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U24 (
    .in(_U24_in),
    .clk(_U24_clk),
    .out(_U24_out)
);
assign _U25_in = _U24_out;
assign _U25_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U25 (
    .in(_U25_in),
    .clk(_U25_clk),
    .out(_U25_out)
);
assign _U26_in = _U25_out;
assign _U26_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U26 (
    .in(_U26_in),
    .clk(_U26_clk),
    .out(_U26_out)
);
assign _U27_in = _U29_out;
_U27_pt__U28 _U27 (
    .in(_U27_in),
    .out(_U27_out)
);
assign _U29_in = 16'(_U33_out + _U45_out);
assign _U29_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U29 (
    .in(_U29_in),
    .clk(_U29_clk),
    .out(_U29_out)
);
assign _U30_in = _U32_out;
_U30_pt__U31 _U30 (
    .in(_U30_in),
    .out(_U30_out)
);
assign _U32_in = 16'(_U13_out + _U27_out);
assign _U32_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U32 (
    .in(_U32_in),
    .clk(_U32_clk),
    .out(_U32_out)
);
assign _U33_in = _U44_out;
_U33_pt__U34 _U33 (
    .in(_U33_in),
    .out(_U33_out)
);
assign _U35_in = 16'(_U107_out * _U110_out);
assign _U35_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U35 (
    .in(_U35_in),
    .clk(_U35_clk),
    .out(_U35_out)
);
assign _U36_in = _U35_out;
assign _U36_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(_U36_in),
    .clk(_U36_clk),
    .out(_U36_out)
);
assign _U37_in = _U36_out;
assign _U37_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U37 (
    .in(_U37_in),
    .clk(_U37_clk),
    .out(_U37_out)
);
assign _U38_in = _U37_out;
assign _U38_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U38 (
    .in(_U38_in),
    .clk(_U38_clk),
    .out(_U38_out)
);
assign _U39_in = _U38_out;
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign _U4_in = _U6_out;
_U4_pt__U5 _U4 (
    .in(_U4_in),
    .out(_U4_out)
);
assign _U40_in = _U39_out;
assign _U40_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U40 (
    .in(_U40_in),
    .clk(_U40_clk),
    .out(_U40_out)
);
assign _U41_in = _U40_out;
assign _U41_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U41 (
    .in(_U41_in),
    .clk(_U41_clk),
    .out(_U41_out)
);
assign _U42_in = _U41_out;
assign _U42_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U42 (
    .in(_U42_in),
    .clk(_U42_clk),
    .out(_U42_out)
);
assign _U43_in = _U42_out;
assign _U43_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U43 (
    .in(_U43_in),
    .clk(_U43_clk),
    .out(_U43_out)
);
assign _U44_in = _U43_out;
assign _U44_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U44 (
    .in(_U44_in),
    .clk(_U44_clk),
    .out(_U44_out)
);
assign _U45_in = _U47_out;
_U45_pt__U46 _U45 (
    .in(_U45_in),
    .out(_U45_out)
);
assign _U47_in = 16'(_U48_out + _U58_out);
assign _U47_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U47 (
    .in(_U47_in),
    .clk(_U47_clk),
    .out(_U47_out)
);
assign _U48_in = _U57_out;
_U48_pt__U49 _U48 (
    .in(_U48_in),
    .out(_U48_out)
);
assign _U50_in = 16'(_U113_out * _U117_out);
assign _U50_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U50 (
    .in(_U50_in),
    .clk(_U50_clk),
    .out(_U50_out)
);
assign _U51_in = _U50_out;
assign _U51_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U51 (
    .in(_U51_in),
    .clk(_U51_clk),
    .out(_U51_out)
);
assign _U52_in = _U51_out;
assign _U52_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U52 (
    .in(_U52_in),
    .clk(_U52_clk),
    .out(_U52_out)
);
assign _U53_in = _U52_out;
assign _U53_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U53 (
    .in(_U53_in),
    .clk(_U53_clk),
    .out(_U53_out)
);
assign _U54_in = _U53_out;
assign _U54_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U54 (
    .in(_U54_in),
    .clk(_U54_clk),
    .out(_U54_out)
);
assign _U55_in = _U54_out;
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign _U56_in = _U55_out;
assign _U56_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U56 (
    .in(_U56_in),
    .clk(_U56_clk),
    .out(_U56_out)
);
assign _U57_in = _U56_out;
assign _U57_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U57 (
    .in(_U57_in),
    .clk(_U57_clk),
    .out(_U57_out)
);
assign _U58_in = _U60_out;
_U58_pt__U59 _U58 (
    .in(_U58_in),
    .out(_U58_out)
);
assign _U6_in = 16'(_U173_out * _U189_out);
assign _U6_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U6 (
    .in(_U6_in),
    .clk(_U6_clk),
    .out(_U6_out)
);
assign _U60_in = 16'(_U61_out + _U69_out);
assign _U60_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U60 (
    .in(_U60_in),
    .clk(_U60_clk),
    .out(_U60_out)
);
assign _U61_in = _U68_out;
_U61_pt__U62 _U61 (
    .in(_U61_in),
    .out(_U61_out)
);
assign _U63_in = 16'(_U121_out * _U126_out);
assign _U63_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U63 (
    .in(_U63_in),
    .clk(_U63_clk),
    .out(_U63_out)
);
assign _U64_in = _U63_out;
assign _U64_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U64 (
    .in(_U64_in),
    .clk(_U64_clk),
    .out(_U64_out)
);
assign _U65_in = _U64_out;
assign _U65_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U65 (
    .in(_U65_in),
    .clk(_U65_clk),
    .out(_U65_out)
);
assign _U66_in = _U65_out;
assign _U66_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(_U66_in),
    .clk(_U66_clk),
    .out(_U66_out)
);
assign _U67_in = _U66_out;
assign _U67_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U67 (
    .in(_U67_in),
    .clk(_U67_clk),
    .out(_U67_out)
);
assign _U68_in = _U67_out;
assign _U68_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U68 (
    .in(_U68_in),
    .clk(_U68_clk),
    .out(_U68_out)
);
assign _U69_in = _U71_out;
_U69_pt__U70 _U69 (
    .in(_U69_in),
    .out(_U69_out)
);
assign _U7_in = _U10_out;
_U7_pt__U8 _U7 (
    .in(_U7_in),
    .out(_U7_out)
);
assign _U71_in = 16'(_U72_out + _U78_out);
assign _U71_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U71 (
    .in(_U71_in),
    .clk(_U71_clk),
    .out(_U71_out)
);
assign _U72_in = _U77_out;
_U72_pt__U73 _U72 (
    .in(_U72_in),
    .out(_U72_out)
);
assign _U74_in = 16'(_U131_out * _U137_out);
assign _U74_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U74 (
    .in(_U74_in),
    .clk(_U74_clk),
    .out(_U74_out)
);
assign _U75_in = _U74_out;
assign _U75_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U75 (
    .in(_U75_in),
    .clk(_U75_clk),
    .out(_U75_out)
);
assign _U76_in = _U75_out;
assign _U76_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U76 (
    .in(_U76_in),
    .clk(_U76_clk),
    .out(_U76_out)
);
assign _U77_in = _U76_out;
assign _U77_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(_U77_in),
    .clk(_U77_clk),
    .out(_U77_out)
);
assign _U78_in = _U80_out;
_U78_pt__U79 _U78 (
    .in(_U78_in),
    .out(_U78_out)
);
assign _U80_in = 16'(_U81_out + _U85_out);
assign _U80_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(_U80_in),
    .clk(_U80_clk),
    .out(_U80_out)
);
assign _U81_in = _U84_out;
_U81_pt__U82 _U81 (
    .in(_U81_in),
    .out(_U81_out)
);
assign _U83_in = 16'(_U143_out * _U150_out);
assign _U83_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U83 (
    .in(_U83_in),
    .clk(_U83_clk),
    .out(_U83_out)
);
assign _U84_in = _U83_out;
assign _U84_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U84 (
    .in(_U84_in),
    .clk(_U84_clk),
    .out(_U84_out)
);
assign _U85_in = _U87_out;
_U85_pt__U86 _U85 (
    .in(_U85_in),
    .out(_U85_out)
);
assign _U87_in = 16'(_U157_out * _U165_out);
assign _U87_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U87 (
    .in(_U87_in),
    .clk(_U87_clk),
    .out(_U87_out)
);
assign _U88_in = _U102_out;
_U88_pt__U89 _U88 (
    .in(_U88_in),
    .out(_U88_out)
);
assign _U9_in = 16'(_U88_out + _U30_out);
assign _U9_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U9 (
    .in(_U9_in),
    .clk(_U9_clk),
    .out(_U9_out)
);
assign _U90_in = in0_conv_stencil[0];
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = _U90_out;
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = _U91_out;
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign _U93_in = _U92_out;
assign _U93_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U93_in),
    .clk(_U93_clk),
    .out(_U93_out)
);
assign _U94_in = _U93_out;
assign _U94_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U94_in),
    .clk(_U94_clk),
    .out(_U94_out)
);
assign _U95_in = _U94_out;
assign _U95_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U95 (
    .in(_U95_in),
    .clk(_U95_clk),
    .out(_U95_out)
);
assign _U96_in = _U95_out;
assign _U96_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U96 (
    .in(_U96_in),
    .clk(_U96_clk),
    .out(_U96_out)
);
assign _U97_in = _U96_out;
assign _U97_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(_U97_in),
    .clk(_U97_clk),
    .out(_U97_out)
);
assign _U98_in = _U97_out;
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = _U98_out;
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U0_pt__U1 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U0_in;
assign _U0_in = in0_hw_input_stencil[0];
_U0_pt__U1 _U0 (
    .in(_U0_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U121_clk;
wire [15:0] arr__U121_in [4:0];
wire [15:0] arr__U121_out [4:0];
wire arr__U128_clk;
wire [15:0] arr__U128_in [4:0];
wire [15:0] arr__U128_out [4:0];
wire arr__U135_clk;
wire [15:0] arr__U135_in [4:0];
wire [15:0] arr__U135_out [4:0];
wire arr__U142_clk;
wire [15:0] arr__U142_in [4:0];
wire [15:0] arr__U142_out [4:0];
wire arr__U149_clk;
wire [15:0] arr__U149_in [4:0];
wire [15:0] arr__U149_out [4:0];
wire arr__U156_clk;
wire [15:0] arr__U156_in [4:0];
wire [15:0] arr__U156_out [4:0];
wire arr__U163_clk;
wire [15:0] arr__U163_in [4:0];
wire [15:0] arr__U163_out [4:0];
wire arr__U170_clk;
wire [15:0] arr__U170_in [4:0];
wire [15:0] arr__U170_out [4:0];
wire arr__U177_clk;
wire [15:0] arr__U177_in [4:0];
wire [15:0] arr__U177_out [4:0];
wire arr__U184_clk;
wire [15:0] arr__U184_in [4:0];
wire [15:0] arr__U184_out [4:0];
wire arr__U191_clk;
wire [15:0] arr__U191_in [4:0];
wire [15:0] arr__U191_out [4:0];
wire arr__U198_clk;
wire [15:0] arr__U198_in [4:0];
wire [15:0] arr__U198_out [4:0];
wire arr__U205_clk;
wire [15:0] arr__U205_in [4:0];
wire [15:0] arr__U205_out [4:0];
wire arr__U212_clk;
wire [15:0] arr__U212_in [4:0];
wire [15:0] arr__U212_out [4:0];
wire arr__U219_clk;
wire [15:0] arr__U219_in [4:0];
wire [15:0] arr__U219_out [4:0];
wire arr__U226_clk;
wire [15:0] arr__U226_in [4:0];
wire [15:0] arr__U226_out [4:0];
wire arr__U233_clk;
wire [15:0] arr__U233_in [4:0];
wire [15:0] arr__U233_out [4:0];
wire arr__U299_clk;
wire [15:0] arr__U299_in [4:0];
wire [15:0] arr__U299_out [4:0];
wire arr__U306_clk;
wire [15:0] arr__U306_in [4:0];
wire [15:0] arr__U306_out [4:0];
wire arr__U332_clk;
wire [15:0] arr__U332_in [4:0];
wire [15:0] arr__U332_out [4:0];
wire arr__U339_clk;
wire [15:0] arr__U339_in [4:0];
wire [15:0] arr__U339_out [4:0];
wire arr__U346_clk;
wire [15:0] arr__U346_in [4:0];
wire [15:0] arr__U346_out [4:0];
wire arr__U353_clk;
wire [15:0] arr__U353_in [4:0];
wire [15:0] arr__U353_out [4:0];
wire arr__U360_clk;
wire [15:0] arr__U360_in [4:0];
wire [15:0] arr__U360_out [4:0];
wire arr__U367_clk;
wire [15:0] arr__U367_in [4:0];
wire [15:0] arr__U367_out [4:0];
wire arr__U374_clk;
wire [15:0] arr__U374_in [4:0];
wire [15:0] arr__U374_out [4:0];
wire arr__U381_clk;
wire [15:0] arr__U381_in [4:0];
wire [15:0] arr__U381_out [4:0];
wire arr__U388_clk;
wire [15:0] arr__U388_in [4:0];
wire [15:0] arr__U388_out [4:0];
wire arr__U395_clk;
wire [15:0] arr__U395_in [4:0];
wire [15:0] arr__U395_out [4:0];
wire arr__U402_clk;
wire [15:0] arr__U402_in [4:0];
wire [15:0] arr__U402_out [4:0];
wire arr__U409_clk;
wire [15:0] arr__U409_in [4:0];
wire [15:0] arr__U409_out [4:0];
wire arr__U416_clk;
wire [15:0] arr__U416_in [4:0];
wire [15:0] arr__U416_out [4:0];
wire arr__U423_clk;
wire [15:0] arr__U423_in [4:0];
wire [15:0] arr__U423_out [4:0];
wire arr__U430_clk;
wire [15:0] arr__U430_in [4:0];
wire [15:0] arr__U430_out [4:0];
wire arr__U437_clk;
wire [15:0] arr__U437_in [4:0];
wire [15:0] arr__U437_out [4:0];
wire arr__U444_clk;
wire [15:0] arr__U444_in [4:0];
wire [15:0] arr__U444_out [4:0];
wire arr__U510_clk;
wire [15:0] arr__U510_in [4:0];
wire [15:0] arr__U510_out [4:0];
wire arr__U517_clk;
wire [15:0] arr__U517_in [4:0];
wire [15:0] arr__U517_out [4:0];
wire arr__U543_clk;
wire [15:0] arr__U543_in [4:0];
wire [15:0] arr__U543_out [4:0];
wire arr__U550_clk;
wire [15:0] arr__U550_in [4:0];
wire [15:0] arr__U550_out [4:0];
wire arr__U557_clk;
wire [15:0] arr__U557_in [4:0];
wire [15:0] arr__U557_out [4:0];
wire arr__U564_clk;
wire [15:0] arr__U564_in [4:0];
wire [15:0] arr__U564_out [4:0];
wire arr__U571_clk;
wire [15:0] arr__U571_in [4:0];
wire [15:0] arr__U571_out [4:0];
wire arr__U578_clk;
wire [15:0] arr__U578_in [4:0];
wire [15:0] arr__U578_out [4:0];
wire arr__U585_clk;
wire [15:0] arr__U585_in [4:0];
wire [15:0] arr__U585_out [4:0];
wire arr__U592_clk;
wire [15:0] arr__U592_in [4:0];
wire [15:0] arr__U592_out [4:0];
wire arr__U599_clk;
wire [15:0] arr__U599_in [4:0];
wire [15:0] arr__U599_out [4:0];
wire arr__U606_clk;
wire [15:0] arr__U606_in [4:0];
wire [15:0] arr__U606_out [4:0];
wire arr__U613_clk;
wire [15:0] arr__U613_in [4:0];
wire [15:0] arr__U613_out [4:0];
wire arr__U620_clk;
wire [15:0] arr__U620_in [4:0];
wire [15:0] arr__U620_out [4:0];
wire arr__U627_clk;
wire [15:0] arr__U627_in [4:0];
wire [15:0] arr__U627_out [4:0];
wire arr__U634_clk;
wire [15:0] arr__U634_in [4:0];
wire [15:0] arr__U634_out [4:0];
wire arr__U641_clk;
wire [15:0] arr__U641_in [4:0];
wire [15:0] arr__U641_out [4:0];
wire arr__U648_clk;
wire [15:0] arr__U648_in [4:0];
wire [15:0] arr__U648_out [4:0];
wire arr__U655_clk;
wire [15:0] arr__U655_in [4:0];
wire [15:0] arr__U655_out [4:0];
wire arr__U727_clk;
wire [15:0] arr__U727_in [3:0];
wire [15:0] arr__U727_out [3:0];
wire arr__U733_clk;
wire [15:0] arr__U733_in [3:0];
wire [15:0] arr__U733_out [3:0];
wire arr__U743_clk;
wire [15:0] arr__U743_in [3:0];
wire [15:0] arr__U743_out [3:0];
wire arr__U749_clk;
wire [15:0] arr__U749_in [3:0];
wire [15:0] arr__U749_out [3:0];
wire arr__U88_clk;
wire [15:0] arr__U88_in [4:0];
wire [15:0] arr__U88_out [4:0];
wire arr__U95_clk;
wire [15:0] arr__U95_in [4:0];
wire [15:0] arr__U95_out [4:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U103_clk;
wire delay_reg__U103_in;
wire delay_reg__U103_out;
wire delay_reg__U104_clk;
wire delay_reg__U104_in;
wire delay_reg__U104_out;
wire delay_reg__U105_clk;
wire delay_reg__U105_in;
wire delay_reg__U105_out;
wire delay_reg__U106_clk;
wire delay_reg__U106_in;
wire delay_reg__U106_out;
wire delay_reg__U107_clk;
wire delay_reg__U107_in;
wire delay_reg__U107_out;
wire delay_reg__U108_clk;
wire delay_reg__U108_in;
wire delay_reg__U108_out;
wire delay_reg__U109_clk;
wire delay_reg__U109_in;
wire delay_reg__U109_out;
wire delay_reg__U110_clk;
wire delay_reg__U110_in;
wire delay_reg__U110_out;
wire delay_reg__U111_clk;
wire delay_reg__U111_in;
wire delay_reg__U111_out;
wire delay_reg__U112_clk;
wire delay_reg__U112_in;
wire delay_reg__U112_out;
wire delay_reg__U113_clk;
wire delay_reg__U113_in;
wire delay_reg__U113_out;
wire delay_reg__U114_clk;
wire delay_reg__U114_in;
wire delay_reg__U114_out;
wire delay_reg__U115_clk;
wire delay_reg__U115_in;
wire delay_reg__U115_out;
wire delay_reg__U116_clk;
wire delay_reg__U116_in;
wire delay_reg__U116_out;
wire delay_reg__U117_clk;
wire delay_reg__U117_in;
wire delay_reg__U117_out;
wire delay_reg__U118_clk;
wire delay_reg__U118_in;
wire delay_reg__U118_out;
wire delay_reg__U119_clk;
wire delay_reg__U119_in;
wire delay_reg__U119_out;
wire delay_reg__U296_clk;
wire delay_reg__U296_in;
wire delay_reg__U296_out;
wire delay_reg__U297_clk;
wire delay_reg__U297_in;
wire delay_reg__U297_out;
wire delay_reg__U314_clk;
wire delay_reg__U314_in;
wire delay_reg__U314_out;
wire delay_reg__U315_clk;
wire delay_reg__U315_in;
wire delay_reg__U315_out;
wire delay_reg__U316_clk;
wire delay_reg__U316_in;
wire delay_reg__U316_out;
wire delay_reg__U317_clk;
wire delay_reg__U317_in;
wire delay_reg__U317_out;
wire delay_reg__U318_clk;
wire delay_reg__U318_in;
wire delay_reg__U318_out;
wire delay_reg__U319_clk;
wire delay_reg__U319_in;
wire delay_reg__U319_out;
wire delay_reg__U320_clk;
wire delay_reg__U320_in;
wire delay_reg__U320_out;
wire delay_reg__U321_clk;
wire delay_reg__U321_in;
wire delay_reg__U321_out;
wire delay_reg__U322_clk;
wire delay_reg__U322_in;
wire delay_reg__U322_out;
wire delay_reg__U323_clk;
wire delay_reg__U323_in;
wire delay_reg__U323_out;
wire delay_reg__U324_clk;
wire delay_reg__U324_in;
wire delay_reg__U324_out;
wire delay_reg__U325_clk;
wire delay_reg__U325_in;
wire delay_reg__U325_out;
wire delay_reg__U326_clk;
wire delay_reg__U326_in;
wire delay_reg__U326_out;
wire delay_reg__U327_clk;
wire delay_reg__U327_in;
wire delay_reg__U327_out;
wire delay_reg__U328_clk;
wire delay_reg__U328_in;
wire delay_reg__U328_out;
wire delay_reg__U329_clk;
wire delay_reg__U329_in;
wire delay_reg__U329_out;
wire delay_reg__U330_clk;
wire delay_reg__U330_in;
wire delay_reg__U330_out;
wire delay_reg__U507_clk;
wire delay_reg__U507_in;
wire delay_reg__U507_out;
wire delay_reg__U508_clk;
wire delay_reg__U508_in;
wire delay_reg__U508_out;
wire delay_reg__U525_clk;
wire delay_reg__U525_in;
wire delay_reg__U525_out;
wire delay_reg__U526_clk;
wire delay_reg__U526_in;
wire delay_reg__U526_out;
wire delay_reg__U527_clk;
wire delay_reg__U527_in;
wire delay_reg__U527_out;
wire delay_reg__U528_clk;
wire delay_reg__U528_in;
wire delay_reg__U528_out;
wire delay_reg__U529_clk;
wire delay_reg__U529_in;
wire delay_reg__U529_out;
wire delay_reg__U530_clk;
wire delay_reg__U530_in;
wire delay_reg__U530_out;
wire delay_reg__U531_clk;
wire delay_reg__U531_in;
wire delay_reg__U531_out;
wire delay_reg__U532_clk;
wire delay_reg__U532_in;
wire delay_reg__U532_out;
wire delay_reg__U533_clk;
wire delay_reg__U533_in;
wire delay_reg__U533_out;
wire delay_reg__U534_clk;
wire delay_reg__U534_in;
wire delay_reg__U534_out;
wire delay_reg__U535_clk;
wire delay_reg__U535_in;
wire delay_reg__U535_out;
wire delay_reg__U536_clk;
wire delay_reg__U536_in;
wire delay_reg__U536_out;
wire delay_reg__U537_clk;
wire delay_reg__U537_in;
wire delay_reg__U537_out;
wire delay_reg__U538_clk;
wire delay_reg__U538_in;
wire delay_reg__U538_out;
wire delay_reg__U539_clk;
wire delay_reg__U539_in;
wire delay_reg__U539_out;
wire delay_reg__U540_clk;
wire delay_reg__U540_in;
wire delay_reg__U540_out;
wire delay_reg__U541_clk;
wire delay_reg__U541_in;
wire delay_reg__U541_out;
wire delay_reg__U724_clk;
wire delay_reg__U724_in;
wire delay_reg__U724_out;
wire delay_reg__U725_clk;
wire delay_reg__U725_in;
wire delay_reg__U725_out;
wire delay_reg__U740_clk;
wire delay_reg__U740_in;
wire delay_reg__U740_out;
wire delay_reg__U741_clk;
wire delay_reg__U741_in;
wire delay_reg__U741_out;
wire delay_reg__U85_clk;
wire delay_reg__U85_in;
wire delay_reg__U85_out;
wire delay_reg__U86_clk;
wire delay_reg__U86_in;
wire delay_reg__U86_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U121_clk = clk;
assign arr__U121_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U121_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U121_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U121_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U121_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U122 arr__U121 (
    .clk(arr__U121_clk),
    .in(arr__U121_in),
    .out(arr__U121_out)
);
assign arr__U128_clk = clk;
assign arr__U128_in[4] = arr__U121_out[4];
assign arr__U128_in[3] = arr__U121_out[3];
assign arr__U128_in[2] = arr__U121_out[2];
assign arr__U128_in[1] = arr__U121_out[1];
assign arr__U128_in[0] = arr__U121_out[0];
array_delay_U129 arr__U128 (
    .clk(arr__U128_clk),
    .in(arr__U128_in),
    .out(arr__U128_out)
);
assign arr__U135_clk = clk;
assign arr__U135_in[4] = arr__U128_out[4];
assign arr__U135_in[3] = arr__U128_out[3];
assign arr__U135_in[2] = arr__U128_out[2];
assign arr__U135_in[1] = arr__U128_out[1];
assign arr__U135_in[0] = arr__U128_out[0];
array_delay_U136 arr__U135 (
    .clk(arr__U135_clk),
    .in(arr__U135_in),
    .out(arr__U135_out)
);
assign arr__U142_clk = clk;
assign arr__U142_in[4] = arr__U135_out[4];
assign arr__U142_in[3] = arr__U135_out[3];
assign arr__U142_in[2] = arr__U135_out[2];
assign arr__U142_in[1] = arr__U135_out[1];
assign arr__U142_in[0] = arr__U135_out[0];
array_delay_U143 arr__U142 (
    .clk(arr__U142_clk),
    .in(arr__U142_in),
    .out(arr__U142_out)
);
assign arr__U149_clk = clk;
assign arr__U149_in[4] = arr__U142_out[4];
assign arr__U149_in[3] = arr__U142_out[3];
assign arr__U149_in[2] = arr__U142_out[2];
assign arr__U149_in[1] = arr__U142_out[1];
assign arr__U149_in[0] = arr__U142_out[0];
array_delay_U150 arr__U149 (
    .clk(arr__U149_clk),
    .in(arr__U149_in),
    .out(arr__U149_out)
);
assign arr__U156_clk = clk;
assign arr__U156_in[4] = arr__U149_out[4];
assign arr__U156_in[3] = arr__U149_out[3];
assign arr__U156_in[2] = arr__U149_out[2];
assign arr__U156_in[1] = arr__U149_out[1];
assign arr__U156_in[0] = arr__U149_out[0];
array_delay_U157 arr__U156 (
    .clk(arr__U156_clk),
    .in(arr__U156_in),
    .out(arr__U156_out)
);
assign arr__U163_clk = clk;
assign arr__U163_in[4] = arr__U156_out[4];
assign arr__U163_in[3] = arr__U156_out[3];
assign arr__U163_in[2] = arr__U156_out[2];
assign arr__U163_in[1] = arr__U156_out[1];
assign arr__U163_in[0] = arr__U156_out[0];
array_delay_U164 arr__U163 (
    .clk(arr__U163_clk),
    .in(arr__U163_in),
    .out(arr__U163_out)
);
assign arr__U170_clk = clk;
assign arr__U170_in[4] = arr__U163_out[4];
assign arr__U170_in[3] = arr__U163_out[3];
assign arr__U170_in[2] = arr__U163_out[2];
assign arr__U170_in[1] = arr__U163_out[1];
assign arr__U170_in[0] = arr__U163_out[0];
array_delay_U171 arr__U170 (
    .clk(arr__U170_clk),
    .in(arr__U170_in),
    .out(arr__U170_out)
);
assign arr__U177_clk = clk;
assign arr__U177_in[4] = arr__U170_out[4];
assign arr__U177_in[3] = arr__U170_out[3];
assign arr__U177_in[2] = arr__U170_out[2];
assign arr__U177_in[1] = arr__U170_out[1];
assign arr__U177_in[0] = arr__U170_out[0];
array_delay_U178 arr__U177 (
    .clk(arr__U177_clk),
    .in(arr__U177_in),
    .out(arr__U177_out)
);
assign arr__U184_clk = clk;
assign arr__U184_in[4] = arr__U177_out[4];
assign arr__U184_in[3] = arr__U177_out[3];
assign arr__U184_in[2] = arr__U177_out[2];
assign arr__U184_in[1] = arr__U177_out[1];
assign arr__U184_in[0] = arr__U177_out[0];
array_delay_U185 arr__U184 (
    .clk(arr__U184_clk),
    .in(arr__U184_in),
    .out(arr__U184_out)
);
assign arr__U191_clk = clk;
assign arr__U191_in[4] = arr__U184_out[4];
assign arr__U191_in[3] = arr__U184_out[3];
assign arr__U191_in[2] = arr__U184_out[2];
assign arr__U191_in[1] = arr__U184_out[1];
assign arr__U191_in[0] = arr__U184_out[0];
array_delay_U192 arr__U191 (
    .clk(arr__U191_clk),
    .in(arr__U191_in),
    .out(arr__U191_out)
);
assign arr__U198_clk = clk;
assign arr__U198_in[4] = arr__U191_out[4];
assign arr__U198_in[3] = arr__U191_out[3];
assign arr__U198_in[2] = arr__U191_out[2];
assign arr__U198_in[1] = arr__U191_out[1];
assign arr__U198_in[0] = arr__U191_out[0];
array_delay_U199 arr__U198 (
    .clk(arr__U198_clk),
    .in(arr__U198_in),
    .out(arr__U198_out)
);
assign arr__U205_clk = clk;
assign arr__U205_in[4] = arr__U198_out[4];
assign arr__U205_in[3] = arr__U198_out[3];
assign arr__U205_in[2] = arr__U198_out[2];
assign arr__U205_in[1] = arr__U198_out[1];
assign arr__U205_in[0] = arr__U198_out[0];
array_delay_U206 arr__U205 (
    .clk(arr__U205_clk),
    .in(arr__U205_in),
    .out(arr__U205_out)
);
assign arr__U212_clk = clk;
assign arr__U212_in[4] = arr__U205_out[4];
assign arr__U212_in[3] = arr__U205_out[3];
assign arr__U212_in[2] = arr__U205_out[2];
assign arr__U212_in[1] = arr__U205_out[1];
assign arr__U212_in[0] = arr__U205_out[0];
array_delay_U213 arr__U212 (
    .clk(arr__U212_clk),
    .in(arr__U212_in),
    .out(arr__U212_out)
);
assign arr__U219_clk = clk;
assign arr__U219_in[4] = arr__U212_out[4];
assign arr__U219_in[3] = arr__U212_out[3];
assign arr__U219_in[2] = arr__U212_out[2];
assign arr__U219_in[1] = arr__U212_out[1];
assign arr__U219_in[0] = arr__U212_out[0];
array_delay_U220 arr__U219 (
    .clk(arr__U219_clk),
    .in(arr__U219_in),
    .out(arr__U219_out)
);
assign arr__U226_clk = clk;
assign arr__U226_in[4] = arr__U219_out[4];
assign arr__U226_in[3] = arr__U219_out[3];
assign arr__U226_in[2] = arr__U219_out[2];
assign arr__U226_in[1] = arr__U219_out[1];
assign arr__U226_in[0] = arr__U219_out[0];
array_delay_U227 arr__U226 (
    .clk(arr__U226_clk),
    .in(arr__U226_in),
    .out(arr__U226_out)
);
assign arr__U233_clk = clk;
assign arr__U233_in[4] = arr__U226_out[4];
assign arr__U233_in[3] = arr__U226_out[3];
assign arr__U233_in[2] = arr__U226_out[2];
assign arr__U233_in[1] = arr__U226_out[1];
assign arr__U233_in[0] = arr__U226_out[0];
array_delay_U234 arr__U233 (
    .clk(arr__U233_clk),
    .in(arr__U233_in),
    .out(arr__U233_out)
);
assign arr__U299_clk = clk;
assign arr__U299_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U299_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U299_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U299_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U299_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U300 arr__U299 (
    .clk(arr__U299_clk),
    .in(arr__U299_in),
    .out(arr__U299_out)
);
assign arr__U306_clk = clk;
assign arr__U306_in[4] = arr__U299_out[4];
assign arr__U306_in[3] = arr__U299_out[3];
assign arr__U306_in[2] = arr__U299_out[2];
assign arr__U306_in[1] = arr__U299_out[1];
assign arr__U306_in[0] = arr__U299_out[0];
array_delay_U307 arr__U306 (
    .clk(arr__U306_clk),
    .in(arr__U306_in),
    .out(arr__U306_out)
);
assign arr__U332_clk = clk;
assign arr__U332_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U332_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U332_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U332_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U332_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U333 arr__U332 (
    .clk(arr__U332_clk),
    .in(arr__U332_in),
    .out(arr__U332_out)
);
assign arr__U339_clk = clk;
assign arr__U339_in[4] = arr__U332_out[4];
assign arr__U339_in[3] = arr__U332_out[3];
assign arr__U339_in[2] = arr__U332_out[2];
assign arr__U339_in[1] = arr__U332_out[1];
assign arr__U339_in[0] = arr__U332_out[0];
array_delay_U340 arr__U339 (
    .clk(arr__U339_clk),
    .in(arr__U339_in),
    .out(arr__U339_out)
);
assign arr__U346_clk = clk;
assign arr__U346_in[4] = arr__U339_out[4];
assign arr__U346_in[3] = arr__U339_out[3];
assign arr__U346_in[2] = arr__U339_out[2];
assign arr__U346_in[1] = arr__U339_out[1];
assign arr__U346_in[0] = arr__U339_out[0];
array_delay_U347 arr__U346 (
    .clk(arr__U346_clk),
    .in(arr__U346_in),
    .out(arr__U346_out)
);
assign arr__U353_clk = clk;
assign arr__U353_in[4] = arr__U346_out[4];
assign arr__U353_in[3] = arr__U346_out[3];
assign arr__U353_in[2] = arr__U346_out[2];
assign arr__U353_in[1] = arr__U346_out[1];
assign arr__U353_in[0] = arr__U346_out[0];
array_delay_U354 arr__U353 (
    .clk(arr__U353_clk),
    .in(arr__U353_in),
    .out(arr__U353_out)
);
assign arr__U360_clk = clk;
assign arr__U360_in[4] = arr__U353_out[4];
assign arr__U360_in[3] = arr__U353_out[3];
assign arr__U360_in[2] = arr__U353_out[2];
assign arr__U360_in[1] = arr__U353_out[1];
assign arr__U360_in[0] = arr__U353_out[0];
array_delay_U361 arr__U360 (
    .clk(arr__U360_clk),
    .in(arr__U360_in),
    .out(arr__U360_out)
);
assign arr__U367_clk = clk;
assign arr__U367_in[4] = arr__U360_out[4];
assign arr__U367_in[3] = arr__U360_out[3];
assign arr__U367_in[2] = arr__U360_out[2];
assign arr__U367_in[1] = arr__U360_out[1];
assign arr__U367_in[0] = arr__U360_out[0];
array_delay_U368 arr__U367 (
    .clk(arr__U367_clk),
    .in(arr__U367_in),
    .out(arr__U367_out)
);
assign arr__U374_clk = clk;
assign arr__U374_in[4] = arr__U367_out[4];
assign arr__U374_in[3] = arr__U367_out[3];
assign arr__U374_in[2] = arr__U367_out[2];
assign arr__U374_in[1] = arr__U367_out[1];
assign arr__U374_in[0] = arr__U367_out[0];
array_delay_U375 arr__U374 (
    .clk(arr__U374_clk),
    .in(arr__U374_in),
    .out(arr__U374_out)
);
assign arr__U381_clk = clk;
assign arr__U381_in[4] = arr__U374_out[4];
assign arr__U381_in[3] = arr__U374_out[3];
assign arr__U381_in[2] = arr__U374_out[2];
assign arr__U381_in[1] = arr__U374_out[1];
assign arr__U381_in[0] = arr__U374_out[0];
array_delay_U382 arr__U381 (
    .clk(arr__U381_clk),
    .in(arr__U381_in),
    .out(arr__U381_out)
);
assign arr__U388_clk = clk;
assign arr__U388_in[4] = arr__U381_out[4];
assign arr__U388_in[3] = arr__U381_out[3];
assign arr__U388_in[2] = arr__U381_out[2];
assign arr__U388_in[1] = arr__U381_out[1];
assign arr__U388_in[0] = arr__U381_out[0];
array_delay_U389 arr__U388 (
    .clk(arr__U388_clk),
    .in(arr__U388_in),
    .out(arr__U388_out)
);
assign arr__U395_clk = clk;
assign arr__U395_in[4] = arr__U388_out[4];
assign arr__U395_in[3] = arr__U388_out[3];
assign arr__U395_in[2] = arr__U388_out[2];
assign arr__U395_in[1] = arr__U388_out[1];
assign arr__U395_in[0] = arr__U388_out[0];
array_delay_U396 arr__U395 (
    .clk(arr__U395_clk),
    .in(arr__U395_in),
    .out(arr__U395_out)
);
assign arr__U402_clk = clk;
assign arr__U402_in[4] = arr__U395_out[4];
assign arr__U402_in[3] = arr__U395_out[3];
assign arr__U402_in[2] = arr__U395_out[2];
assign arr__U402_in[1] = arr__U395_out[1];
assign arr__U402_in[0] = arr__U395_out[0];
array_delay_U403 arr__U402 (
    .clk(arr__U402_clk),
    .in(arr__U402_in),
    .out(arr__U402_out)
);
assign arr__U409_clk = clk;
assign arr__U409_in[4] = arr__U402_out[4];
assign arr__U409_in[3] = arr__U402_out[3];
assign arr__U409_in[2] = arr__U402_out[2];
assign arr__U409_in[1] = arr__U402_out[1];
assign arr__U409_in[0] = arr__U402_out[0];
array_delay_U410 arr__U409 (
    .clk(arr__U409_clk),
    .in(arr__U409_in),
    .out(arr__U409_out)
);
assign arr__U416_clk = clk;
assign arr__U416_in[4] = arr__U409_out[4];
assign arr__U416_in[3] = arr__U409_out[3];
assign arr__U416_in[2] = arr__U409_out[2];
assign arr__U416_in[1] = arr__U409_out[1];
assign arr__U416_in[0] = arr__U409_out[0];
array_delay_U417 arr__U416 (
    .clk(arr__U416_clk),
    .in(arr__U416_in),
    .out(arr__U416_out)
);
assign arr__U423_clk = clk;
assign arr__U423_in[4] = arr__U416_out[4];
assign arr__U423_in[3] = arr__U416_out[3];
assign arr__U423_in[2] = arr__U416_out[2];
assign arr__U423_in[1] = arr__U416_out[1];
assign arr__U423_in[0] = arr__U416_out[0];
array_delay_U424 arr__U423 (
    .clk(arr__U423_clk),
    .in(arr__U423_in),
    .out(arr__U423_out)
);
assign arr__U430_clk = clk;
assign arr__U430_in[4] = arr__U423_out[4];
assign arr__U430_in[3] = arr__U423_out[3];
assign arr__U430_in[2] = arr__U423_out[2];
assign arr__U430_in[1] = arr__U423_out[1];
assign arr__U430_in[0] = arr__U423_out[0];
array_delay_U431 arr__U430 (
    .clk(arr__U430_clk),
    .in(arr__U430_in),
    .out(arr__U430_out)
);
assign arr__U437_clk = clk;
assign arr__U437_in[4] = arr__U430_out[4];
assign arr__U437_in[3] = arr__U430_out[3];
assign arr__U437_in[2] = arr__U430_out[2];
assign arr__U437_in[1] = arr__U430_out[1];
assign arr__U437_in[0] = arr__U430_out[0];
array_delay_U438 arr__U437 (
    .clk(arr__U437_clk),
    .in(arr__U437_in),
    .out(arr__U437_out)
);
assign arr__U444_clk = clk;
assign arr__U444_in[4] = arr__U437_out[4];
assign arr__U444_in[3] = arr__U437_out[3];
assign arr__U444_in[2] = arr__U437_out[2];
assign arr__U444_in[1] = arr__U437_out[1];
assign arr__U444_in[0] = arr__U437_out[0];
array_delay_U445 arr__U444 (
    .clk(arr__U444_clk),
    .in(arr__U444_in),
    .out(arr__U444_out)
);
assign arr__U510_clk = clk;
assign arr__U510_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U510_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U510_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U510_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U510_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U511 arr__U510 (
    .clk(arr__U510_clk),
    .in(arr__U510_in),
    .out(arr__U510_out)
);
assign arr__U517_clk = clk;
assign arr__U517_in[4] = arr__U510_out[4];
assign arr__U517_in[3] = arr__U510_out[3];
assign arr__U517_in[2] = arr__U510_out[2];
assign arr__U517_in[1] = arr__U510_out[1];
assign arr__U517_in[0] = arr__U510_out[0];
array_delay_U518 arr__U517 (
    .clk(arr__U517_clk),
    .in(arr__U517_in),
    .out(arr__U517_out)
);
assign arr__U543_clk = clk;
assign arr__U543_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U543_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U543_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U543_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U543_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U544 arr__U543 (
    .clk(arr__U543_clk),
    .in(arr__U543_in),
    .out(arr__U543_out)
);
assign arr__U550_clk = clk;
assign arr__U550_in[4] = arr__U543_out[4];
assign arr__U550_in[3] = arr__U543_out[3];
assign arr__U550_in[2] = arr__U543_out[2];
assign arr__U550_in[1] = arr__U543_out[1];
assign arr__U550_in[0] = arr__U543_out[0];
array_delay_U551 arr__U550 (
    .clk(arr__U550_clk),
    .in(arr__U550_in),
    .out(arr__U550_out)
);
assign arr__U557_clk = clk;
assign arr__U557_in[4] = arr__U550_out[4];
assign arr__U557_in[3] = arr__U550_out[3];
assign arr__U557_in[2] = arr__U550_out[2];
assign arr__U557_in[1] = arr__U550_out[1];
assign arr__U557_in[0] = arr__U550_out[0];
array_delay_U558 arr__U557 (
    .clk(arr__U557_clk),
    .in(arr__U557_in),
    .out(arr__U557_out)
);
assign arr__U564_clk = clk;
assign arr__U564_in[4] = arr__U557_out[4];
assign arr__U564_in[3] = arr__U557_out[3];
assign arr__U564_in[2] = arr__U557_out[2];
assign arr__U564_in[1] = arr__U557_out[1];
assign arr__U564_in[0] = arr__U557_out[0];
array_delay_U565 arr__U564 (
    .clk(arr__U564_clk),
    .in(arr__U564_in),
    .out(arr__U564_out)
);
assign arr__U571_clk = clk;
assign arr__U571_in[4] = arr__U564_out[4];
assign arr__U571_in[3] = arr__U564_out[3];
assign arr__U571_in[2] = arr__U564_out[2];
assign arr__U571_in[1] = arr__U564_out[1];
assign arr__U571_in[0] = arr__U564_out[0];
array_delay_U572 arr__U571 (
    .clk(arr__U571_clk),
    .in(arr__U571_in),
    .out(arr__U571_out)
);
assign arr__U578_clk = clk;
assign arr__U578_in[4] = arr__U571_out[4];
assign arr__U578_in[3] = arr__U571_out[3];
assign arr__U578_in[2] = arr__U571_out[2];
assign arr__U578_in[1] = arr__U571_out[1];
assign arr__U578_in[0] = arr__U571_out[0];
array_delay_U579 arr__U578 (
    .clk(arr__U578_clk),
    .in(arr__U578_in),
    .out(arr__U578_out)
);
assign arr__U585_clk = clk;
assign arr__U585_in[4] = arr__U578_out[4];
assign arr__U585_in[3] = arr__U578_out[3];
assign arr__U585_in[2] = arr__U578_out[2];
assign arr__U585_in[1] = arr__U578_out[1];
assign arr__U585_in[0] = arr__U578_out[0];
array_delay_U586 arr__U585 (
    .clk(arr__U585_clk),
    .in(arr__U585_in),
    .out(arr__U585_out)
);
assign arr__U592_clk = clk;
assign arr__U592_in[4] = arr__U585_out[4];
assign arr__U592_in[3] = arr__U585_out[3];
assign arr__U592_in[2] = arr__U585_out[2];
assign arr__U592_in[1] = arr__U585_out[1];
assign arr__U592_in[0] = arr__U585_out[0];
array_delay_U593 arr__U592 (
    .clk(arr__U592_clk),
    .in(arr__U592_in),
    .out(arr__U592_out)
);
assign arr__U599_clk = clk;
assign arr__U599_in[4] = arr__U592_out[4];
assign arr__U599_in[3] = arr__U592_out[3];
assign arr__U599_in[2] = arr__U592_out[2];
assign arr__U599_in[1] = arr__U592_out[1];
assign arr__U599_in[0] = arr__U592_out[0];
array_delay_U600 arr__U599 (
    .clk(arr__U599_clk),
    .in(arr__U599_in),
    .out(arr__U599_out)
);
assign arr__U606_clk = clk;
assign arr__U606_in[4] = arr__U599_out[4];
assign arr__U606_in[3] = arr__U599_out[3];
assign arr__U606_in[2] = arr__U599_out[2];
assign arr__U606_in[1] = arr__U599_out[1];
assign arr__U606_in[0] = arr__U599_out[0];
array_delay_U607 arr__U606 (
    .clk(arr__U606_clk),
    .in(arr__U606_in),
    .out(arr__U606_out)
);
assign arr__U613_clk = clk;
assign arr__U613_in[4] = arr__U606_out[4];
assign arr__U613_in[3] = arr__U606_out[3];
assign arr__U613_in[2] = arr__U606_out[2];
assign arr__U613_in[1] = arr__U606_out[1];
assign arr__U613_in[0] = arr__U606_out[0];
array_delay_U614 arr__U613 (
    .clk(arr__U613_clk),
    .in(arr__U613_in),
    .out(arr__U613_out)
);
assign arr__U620_clk = clk;
assign arr__U620_in[4] = arr__U613_out[4];
assign arr__U620_in[3] = arr__U613_out[3];
assign arr__U620_in[2] = arr__U613_out[2];
assign arr__U620_in[1] = arr__U613_out[1];
assign arr__U620_in[0] = arr__U613_out[0];
array_delay_U621 arr__U620 (
    .clk(arr__U620_clk),
    .in(arr__U620_in),
    .out(arr__U620_out)
);
assign arr__U627_clk = clk;
assign arr__U627_in[4] = arr__U620_out[4];
assign arr__U627_in[3] = arr__U620_out[3];
assign arr__U627_in[2] = arr__U620_out[2];
assign arr__U627_in[1] = arr__U620_out[1];
assign arr__U627_in[0] = arr__U620_out[0];
array_delay_U628 arr__U627 (
    .clk(arr__U627_clk),
    .in(arr__U627_in),
    .out(arr__U627_out)
);
assign arr__U634_clk = clk;
assign arr__U634_in[4] = arr__U627_out[4];
assign arr__U634_in[3] = arr__U627_out[3];
assign arr__U634_in[2] = arr__U627_out[2];
assign arr__U634_in[1] = arr__U627_out[1];
assign arr__U634_in[0] = arr__U627_out[0];
array_delay_U635 arr__U634 (
    .clk(arr__U634_clk),
    .in(arr__U634_in),
    .out(arr__U634_out)
);
assign arr__U641_clk = clk;
assign arr__U641_in[4] = arr__U634_out[4];
assign arr__U641_in[3] = arr__U634_out[3];
assign arr__U641_in[2] = arr__U634_out[2];
assign arr__U641_in[1] = arr__U634_out[1];
assign arr__U641_in[0] = arr__U634_out[0];
array_delay_U642 arr__U641 (
    .clk(arr__U641_clk),
    .in(arr__U641_in),
    .out(arr__U641_out)
);
assign arr__U648_clk = clk;
assign arr__U648_in[4] = arr__U641_out[4];
assign arr__U648_in[3] = arr__U641_out[3];
assign arr__U648_in[2] = arr__U641_out[2];
assign arr__U648_in[1] = arr__U641_out[1];
assign arr__U648_in[0] = arr__U641_out[0];
array_delay_U649 arr__U648 (
    .clk(arr__U648_clk),
    .in(arr__U648_in),
    .out(arr__U648_out)
);
assign arr__U655_clk = clk;
assign arr__U655_in[4] = arr__U648_out[4];
assign arr__U655_in[3] = arr__U648_out[3];
assign arr__U655_in[2] = arr__U648_out[2];
assign arr__U655_in[1] = arr__U648_out[1];
assign arr__U655_in[0] = arr__U648_out[0];
array_delay_U656 arr__U655 (
    .clk(arr__U655_clk),
    .in(arr__U655_in),
    .out(arr__U655_out)
);
assign arr__U727_clk = clk;
assign arr__U727_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U727_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U727_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U727_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U728 arr__U727 (
    .clk(arr__U727_clk),
    .in(arr__U727_in),
    .out(arr__U727_out)
);
assign arr__U733_clk = clk;
assign arr__U733_in[3] = arr__U727_out[3];
assign arr__U733_in[2] = arr__U727_out[2];
assign arr__U733_in[1] = arr__U727_out[1];
assign arr__U733_in[0] = arr__U727_out[0];
array_delay_U734 arr__U733 (
    .clk(arr__U733_clk),
    .in(arr__U733_in),
    .out(arr__U733_out)
);
assign arr__U743_clk = clk;
assign arr__U743_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U743_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U743_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U743_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U744 arr__U743 (
    .clk(arr__U743_clk),
    .in(arr__U743_in),
    .out(arr__U743_out)
);
assign arr__U749_clk = clk;
assign arr__U749_in[3] = arr__U743_out[3];
assign arr__U749_in[2] = arr__U743_out[2];
assign arr__U749_in[1] = arr__U743_out[1];
assign arr__U749_in[0] = arr__U743_out[0];
array_delay_U750 arr__U749 (
    .clk(arr__U749_clk),
    .in(arr__U749_in),
    .out(arr__U749_out)
);
assign arr__U88_clk = clk;
assign arr__U88_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U88_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U88_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U88_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U88_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U89 arr__U88 (
    .clk(arr__U88_clk),
    .in(arr__U88_in),
    .out(arr__U88_out)
);
assign arr__U95_clk = clk;
assign arr__U95_in[4] = arr__U88_out[4];
assign arr__U95_in[3] = arr__U88_out[3];
assign arr__U95_in[2] = arr__U88_out[2];
assign arr__U95_in[1] = arr__U88_out[1];
assign arr__U95_in[0] = arr__U88_out[0];
array_delay_U96 arr__U95 (
    .clk(arr__U95_clk),
    .in(arr__U95_in),
    .out(arr__U95_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U103_clk = clk;
assign delay_reg__U103_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U103 (
    .clk(delay_reg__U103_clk),
    .in(delay_reg__U103_in),
    .out(delay_reg__U103_out)
);
assign delay_reg__U104_clk = clk;
assign delay_reg__U104_in = delay_reg__U103_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U104 (
    .clk(delay_reg__U104_clk),
    .in(delay_reg__U104_in),
    .out(delay_reg__U104_out)
);
assign delay_reg__U105_clk = clk;
assign delay_reg__U105_in = delay_reg__U104_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U105 (
    .clk(delay_reg__U105_clk),
    .in(delay_reg__U105_in),
    .out(delay_reg__U105_out)
);
assign delay_reg__U106_clk = clk;
assign delay_reg__U106_in = delay_reg__U105_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U106 (
    .clk(delay_reg__U106_clk),
    .in(delay_reg__U106_in),
    .out(delay_reg__U106_out)
);
assign delay_reg__U107_clk = clk;
assign delay_reg__U107_in = delay_reg__U106_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U107 (
    .clk(delay_reg__U107_clk),
    .in(delay_reg__U107_in),
    .out(delay_reg__U107_out)
);
assign delay_reg__U108_clk = clk;
assign delay_reg__U108_in = delay_reg__U107_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U108 (
    .clk(delay_reg__U108_clk),
    .in(delay_reg__U108_in),
    .out(delay_reg__U108_out)
);
assign delay_reg__U109_clk = clk;
assign delay_reg__U109_in = delay_reg__U108_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U109 (
    .clk(delay_reg__U109_clk),
    .in(delay_reg__U109_in),
    .out(delay_reg__U109_out)
);
assign delay_reg__U110_clk = clk;
assign delay_reg__U110_in = delay_reg__U109_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U110 (
    .clk(delay_reg__U110_clk),
    .in(delay_reg__U110_in),
    .out(delay_reg__U110_out)
);
assign delay_reg__U111_clk = clk;
assign delay_reg__U111_in = delay_reg__U110_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U111 (
    .clk(delay_reg__U111_clk),
    .in(delay_reg__U111_in),
    .out(delay_reg__U111_out)
);
assign delay_reg__U112_clk = clk;
assign delay_reg__U112_in = delay_reg__U111_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U112 (
    .clk(delay_reg__U112_clk),
    .in(delay_reg__U112_in),
    .out(delay_reg__U112_out)
);
assign delay_reg__U113_clk = clk;
assign delay_reg__U113_in = delay_reg__U112_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U113 (
    .clk(delay_reg__U113_clk),
    .in(delay_reg__U113_in),
    .out(delay_reg__U113_out)
);
assign delay_reg__U114_clk = clk;
assign delay_reg__U114_in = delay_reg__U113_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U114 (
    .clk(delay_reg__U114_clk),
    .in(delay_reg__U114_in),
    .out(delay_reg__U114_out)
);
assign delay_reg__U115_clk = clk;
assign delay_reg__U115_in = delay_reg__U114_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U115 (
    .clk(delay_reg__U115_clk),
    .in(delay_reg__U115_in),
    .out(delay_reg__U115_out)
);
assign delay_reg__U116_clk = clk;
assign delay_reg__U116_in = delay_reg__U115_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U116 (
    .clk(delay_reg__U116_clk),
    .in(delay_reg__U116_in),
    .out(delay_reg__U116_out)
);
assign delay_reg__U117_clk = clk;
assign delay_reg__U117_in = delay_reg__U116_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U117 (
    .clk(delay_reg__U117_clk),
    .in(delay_reg__U117_in),
    .out(delay_reg__U117_out)
);
assign delay_reg__U118_clk = clk;
assign delay_reg__U118_in = delay_reg__U117_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U118 (
    .clk(delay_reg__U118_clk),
    .in(delay_reg__U118_in),
    .out(delay_reg__U118_out)
);
assign delay_reg__U119_clk = clk;
assign delay_reg__U119_in = delay_reg__U118_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U119 (
    .clk(delay_reg__U119_clk),
    .in(delay_reg__U119_in),
    .out(delay_reg__U119_out)
);
assign delay_reg__U296_clk = clk;
assign delay_reg__U296_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U296 (
    .clk(delay_reg__U296_clk),
    .in(delay_reg__U296_in),
    .out(delay_reg__U296_out)
);
assign delay_reg__U297_clk = clk;
assign delay_reg__U297_in = delay_reg__U296_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U297 (
    .clk(delay_reg__U297_clk),
    .in(delay_reg__U297_in),
    .out(delay_reg__U297_out)
);
assign delay_reg__U314_clk = clk;
assign delay_reg__U314_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U314 (
    .clk(delay_reg__U314_clk),
    .in(delay_reg__U314_in),
    .out(delay_reg__U314_out)
);
assign delay_reg__U315_clk = clk;
assign delay_reg__U315_in = delay_reg__U314_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U315 (
    .clk(delay_reg__U315_clk),
    .in(delay_reg__U315_in),
    .out(delay_reg__U315_out)
);
assign delay_reg__U316_clk = clk;
assign delay_reg__U316_in = delay_reg__U315_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U316 (
    .clk(delay_reg__U316_clk),
    .in(delay_reg__U316_in),
    .out(delay_reg__U316_out)
);
assign delay_reg__U317_clk = clk;
assign delay_reg__U317_in = delay_reg__U316_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U317 (
    .clk(delay_reg__U317_clk),
    .in(delay_reg__U317_in),
    .out(delay_reg__U317_out)
);
assign delay_reg__U318_clk = clk;
assign delay_reg__U318_in = delay_reg__U317_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U318 (
    .clk(delay_reg__U318_clk),
    .in(delay_reg__U318_in),
    .out(delay_reg__U318_out)
);
assign delay_reg__U319_clk = clk;
assign delay_reg__U319_in = delay_reg__U318_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U319 (
    .clk(delay_reg__U319_clk),
    .in(delay_reg__U319_in),
    .out(delay_reg__U319_out)
);
assign delay_reg__U320_clk = clk;
assign delay_reg__U320_in = delay_reg__U319_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U320 (
    .clk(delay_reg__U320_clk),
    .in(delay_reg__U320_in),
    .out(delay_reg__U320_out)
);
assign delay_reg__U321_clk = clk;
assign delay_reg__U321_in = delay_reg__U320_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U321 (
    .clk(delay_reg__U321_clk),
    .in(delay_reg__U321_in),
    .out(delay_reg__U321_out)
);
assign delay_reg__U322_clk = clk;
assign delay_reg__U322_in = delay_reg__U321_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U322 (
    .clk(delay_reg__U322_clk),
    .in(delay_reg__U322_in),
    .out(delay_reg__U322_out)
);
assign delay_reg__U323_clk = clk;
assign delay_reg__U323_in = delay_reg__U322_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U323 (
    .clk(delay_reg__U323_clk),
    .in(delay_reg__U323_in),
    .out(delay_reg__U323_out)
);
assign delay_reg__U324_clk = clk;
assign delay_reg__U324_in = delay_reg__U323_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U324 (
    .clk(delay_reg__U324_clk),
    .in(delay_reg__U324_in),
    .out(delay_reg__U324_out)
);
assign delay_reg__U325_clk = clk;
assign delay_reg__U325_in = delay_reg__U324_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U325 (
    .clk(delay_reg__U325_clk),
    .in(delay_reg__U325_in),
    .out(delay_reg__U325_out)
);
assign delay_reg__U326_clk = clk;
assign delay_reg__U326_in = delay_reg__U325_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U326 (
    .clk(delay_reg__U326_clk),
    .in(delay_reg__U326_in),
    .out(delay_reg__U326_out)
);
assign delay_reg__U327_clk = clk;
assign delay_reg__U327_in = delay_reg__U326_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U327 (
    .clk(delay_reg__U327_clk),
    .in(delay_reg__U327_in),
    .out(delay_reg__U327_out)
);
assign delay_reg__U328_clk = clk;
assign delay_reg__U328_in = delay_reg__U327_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U328 (
    .clk(delay_reg__U328_clk),
    .in(delay_reg__U328_in),
    .out(delay_reg__U328_out)
);
assign delay_reg__U329_clk = clk;
assign delay_reg__U329_in = delay_reg__U328_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U329 (
    .clk(delay_reg__U329_clk),
    .in(delay_reg__U329_in),
    .out(delay_reg__U329_out)
);
assign delay_reg__U330_clk = clk;
assign delay_reg__U330_in = delay_reg__U329_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U330 (
    .clk(delay_reg__U330_clk),
    .in(delay_reg__U330_in),
    .out(delay_reg__U330_out)
);
assign delay_reg__U507_clk = clk;
assign delay_reg__U507_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U507 (
    .clk(delay_reg__U507_clk),
    .in(delay_reg__U507_in),
    .out(delay_reg__U507_out)
);
assign delay_reg__U508_clk = clk;
assign delay_reg__U508_in = delay_reg__U507_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U508 (
    .clk(delay_reg__U508_clk),
    .in(delay_reg__U508_in),
    .out(delay_reg__U508_out)
);
assign delay_reg__U525_clk = clk;
assign delay_reg__U525_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U525 (
    .clk(delay_reg__U525_clk),
    .in(delay_reg__U525_in),
    .out(delay_reg__U525_out)
);
assign delay_reg__U526_clk = clk;
assign delay_reg__U526_in = delay_reg__U525_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U526 (
    .clk(delay_reg__U526_clk),
    .in(delay_reg__U526_in),
    .out(delay_reg__U526_out)
);
assign delay_reg__U527_clk = clk;
assign delay_reg__U527_in = delay_reg__U526_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U527 (
    .clk(delay_reg__U527_clk),
    .in(delay_reg__U527_in),
    .out(delay_reg__U527_out)
);
assign delay_reg__U528_clk = clk;
assign delay_reg__U528_in = delay_reg__U527_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U528 (
    .clk(delay_reg__U528_clk),
    .in(delay_reg__U528_in),
    .out(delay_reg__U528_out)
);
assign delay_reg__U529_clk = clk;
assign delay_reg__U529_in = delay_reg__U528_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U529 (
    .clk(delay_reg__U529_clk),
    .in(delay_reg__U529_in),
    .out(delay_reg__U529_out)
);
assign delay_reg__U530_clk = clk;
assign delay_reg__U530_in = delay_reg__U529_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U530 (
    .clk(delay_reg__U530_clk),
    .in(delay_reg__U530_in),
    .out(delay_reg__U530_out)
);
assign delay_reg__U531_clk = clk;
assign delay_reg__U531_in = delay_reg__U530_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U531 (
    .clk(delay_reg__U531_clk),
    .in(delay_reg__U531_in),
    .out(delay_reg__U531_out)
);
assign delay_reg__U532_clk = clk;
assign delay_reg__U532_in = delay_reg__U531_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U532 (
    .clk(delay_reg__U532_clk),
    .in(delay_reg__U532_in),
    .out(delay_reg__U532_out)
);
assign delay_reg__U533_clk = clk;
assign delay_reg__U533_in = delay_reg__U532_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U533 (
    .clk(delay_reg__U533_clk),
    .in(delay_reg__U533_in),
    .out(delay_reg__U533_out)
);
assign delay_reg__U534_clk = clk;
assign delay_reg__U534_in = delay_reg__U533_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U534 (
    .clk(delay_reg__U534_clk),
    .in(delay_reg__U534_in),
    .out(delay_reg__U534_out)
);
assign delay_reg__U535_clk = clk;
assign delay_reg__U535_in = delay_reg__U534_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U535 (
    .clk(delay_reg__U535_clk),
    .in(delay_reg__U535_in),
    .out(delay_reg__U535_out)
);
assign delay_reg__U536_clk = clk;
assign delay_reg__U536_in = delay_reg__U535_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U536 (
    .clk(delay_reg__U536_clk),
    .in(delay_reg__U536_in),
    .out(delay_reg__U536_out)
);
assign delay_reg__U537_clk = clk;
assign delay_reg__U537_in = delay_reg__U536_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U537 (
    .clk(delay_reg__U537_clk),
    .in(delay_reg__U537_in),
    .out(delay_reg__U537_out)
);
assign delay_reg__U538_clk = clk;
assign delay_reg__U538_in = delay_reg__U537_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U538 (
    .clk(delay_reg__U538_clk),
    .in(delay_reg__U538_in),
    .out(delay_reg__U538_out)
);
assign delay_reg__U539_clk = clk;
assign delay_reg__U539_in = delay_reg__U538_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U539 (
    .clk(delay_reg__U539_clk),
    .in(delay_reg__U539_in),
    .out(delay_reg__U539_out)
);
assign delay_reg__U540_clk = clk;
assign delay_reg__U540_in = delay_reg__U539_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U540 (
    .clk(delay_reg__U540_clk),
    .in(delay_reg__U540_in),
    .out(delay_reg__U540_out)
);
assign delay_reg__U541_clk = clk;
assign delay_reg__U541_in = delay_reg__U540_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U541 (
    .clk(delay_reg__U541_clk),
    .in(delay_reg__U541_in),
    .out(delay_reg__U541_out)
);
assign delay_reg__U724_clk = clk;
assign delay_reg__U724_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U724 (
    .clk(delay_reg__U724_clk),
    .in(delay_reg__U724_in),
    .out(delay_reg__U724_out)
);
assign delay_reg__U725_clk = clk;
assign delay_reg__U725_in = delay_reg__U724_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U725 (
    .clk(delay_reg__U725_clk),
    .in(delay_reg__U725_in),
    .out(delay_reg__U725_out)
);
assign delay_reg__U740_clk = clk;
assign delay_reg__U740_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U740 (
    .clk(delay_reg__U740_clk),
    .in(delay_reg__U740_in),
    .out(delay_reg__U740_out)
);
assign delay_reg__U741_clk = clk;
assign delay_reg__U741_in = delay_reg__U740_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U741 (
    .clk(delay_reg__U741_clk),
    .in(delay_reg__U741_in),
    .out(delay_reg__U741_out)
);
assign delay_reg__U85_clk = clk;
assign delay_reg__U85_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U85 (
    .clk(delay_reg__U85_clk),
    .in(delay_reg__U85_in),
    .out(delay_reg__U85_out)
);
assign delay_reg__U86_clk = clk;
assign delay_reg__U86_in = delay_reg__U85_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U86 (
    .clk(delay_reg__U86_clk),
    .in(delay_reg__U86_in),
    .out(delay_reg__U86_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U48 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U49 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
affine_controller__U29 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U46 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U47 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U50 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U51 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U470 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U471 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
affine_controller__U451 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U468 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U469 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U472 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U473 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U508_out;
op_hcompute_conv_stencil_3_exe_start_pt__U506 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U517_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U517_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U517_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U517_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U517_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U509 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
affine_controller__U474 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U504 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U505 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U541_out;
op_hcompute_conv_stencil_3_write_start_pt__U524 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U655_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U655_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U655_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U655_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U655_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U542 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U86_out;
op_hcompute_conv_stencil_4_exe_start_pt__U84 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U95_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U95_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U95_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U95_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U95_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U87 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
affine_controller__U52 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U82 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U83 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U119_out;
op_hcompute_conv_stencil_4_write_start_pt__U102 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U233_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U233_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U233_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U233_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U233_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U120 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U297_out;
op_hcompute_conv_stencil_5_exe_start_pt__U295 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U306_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U306_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U306_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U306_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U306_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U298 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
affine_controller__U263 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U293 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U294 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U330_out;
op_hcompute_conv_stencil_5_write_start_pt__U313 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U444_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U444_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U444_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U444_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U444_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U331 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U259 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U260 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
affine_controller__U240 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U257 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U258 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U261 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U262 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U25 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U26 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U0 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U23 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U24 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U27 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U28 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U694 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U695 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U662 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U692 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U693 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U696 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U697 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U725_out;
op_hcompute_hw_output_stencil_exe_start_pt__U723 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U733_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U733_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U733_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U733_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U726 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
affine_controller__U698 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U721 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U722 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U741_out;
op_hcompute_hw_output_stencil_write_start_pt__U739 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U749_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U749_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U749_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U749_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U742 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

