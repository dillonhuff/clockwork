// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
// Module `affine_controller__U88` defined externally
// Module `affine_controller__U81` defined externally
// Module `affine_controller__U7` defined externally
// Module `affine_controller__U60` defined externally
// Module `affine_controller__U37` defined externally
// Module `affine_controller__U14` defined externally
// Module `affine_controller__U118` defined externally
// Module `affine_controller__U111` defined externally
// Module `affine_controller__U0` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U72 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U74 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U61 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U62 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U63 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U65 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U116 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U117 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U112 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U113 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U114 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U115 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U86 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U87 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U82 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U83 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U84 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U85 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U123 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U124 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U119 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U120 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U121 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U122 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U50 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U52 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U38 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U39 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U42 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U27 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U29 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U15 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U16 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U17 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U19 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U101 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U103 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U89 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U90 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U91 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U93 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U12 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U13 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U8 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U9 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U10 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U11 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U5 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U6 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U1 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U2 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U3 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U4 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module hcompute_hw_output_stencil (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
assign out_hw_output_stencil = in0_conv_stencil[0];
endmodule

module hcompute_hw_kernel_global_wrapper_stencil (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
assign out_hw_kernel_global_wrapper_stencil = in0_hw_kernel_stencil[0];
endmodule

module hcompute_hw_input_global_wrapper_stencil (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
assign out_hw_input_global_wrapper_stencil = in0_hw_input_stencil[0];
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module hcompute_conv_stencil_2 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_1 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_5 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_4 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_3 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U95 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U96_in;
wire _U96_clk;
wire [15:0] _U96_out;
wire [15:0] _U97_in;
wire _U97_clk;
wire [15:0] _U97_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U100_in = in[4];
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U96_in = in[0];
assign _U96_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U96 (
    .in(_U96_in),
    .clk(_U96_clk),
    .out(_U96_out)
);
assign _U97_in = in[1];
assign _U97_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(_U97_in),
    .clk(_U97_clk),
    .out(_U97_out)
);
assign _U98_in = in[2];
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = in[3];
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
assign out[4] = _U100_out;
assign out[3] = _U99_out;
assign out[2] = _U98_out;
assign out[1] = _U97_out;
assign out[0] = _U96_out;
endmodule

module array_delay_U76 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U77_in;
wire _U77_clk;
wire [15:0] _U77_out;
wire [15:0] _U78_in;
wire _U78_clk;
wire [15:0] _U78_out;
wire [15:0] _U79_in;
wire _U79_clk;
wire [15:0] _U79_out;
wire [15:0] _U80_in;
wire _U80_clk;
wire [15:0] _U80_out;
assign _U77_in = in[0];
assign _U77_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(_U77_in),
    .clk(_U77_clk),
    .out(_U77_out)
);
assign _U78_in = in[1];
assign _U78_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U78 (
    .in(_U78_in),
    .clk(_U78_clk),
    .out(_U78_out)
);
assign _U79_in = in[2];
assign _U79_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(_U79_in),
    .clk(_U79_clk),
    .out(_U79_out)
);
assign _U80_in = in[3];
assign _U80_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(_U80_in),
    .clk(_U80_clk),
    .out(_U80_out)
);
assign out[3] = _U80_out;
assign out[2] = _U79_out;
assign out[1] = _U78_out;
assign out[0] = _U77_out;
endmodule

module array_delay_U67 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U68_in;
wire _U68_clk;
wire [15:0] _U68_out;
wire [15:0] _U69_in;
wire _U69_clk;
wire [15:0] _U69_out;
wire [15:0] _U70_in;
wire _U70_clk;
wire [15:0] _U70_out;
wire [15:0] _U71_in;
wire _U71_clk;
wire [15:0] _U71_out;
assign _U68_in = in[0];
assign _U68_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U68 (
    .in(_U68_in),
    .clk(_U68_clk),
    .out(_U68_out)
);
assign _U69_in = in[1];
assign _U69_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(_U69_in),
    .clk(_U69_clk),
    .out(_U69_out)
);
assign _U70_in = in[2];
assign _U70_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U70 (
    .in(_U70_in),
    .clk(_U70_clk),
    .out(_U70_out)
);
assign _U71_in = in[3];
assign _U71_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U71 (
    .in(_U71_in),
    .clk(_U71_clk),
    .out(_U71_out)
);
assign out[3] = _U71_out;
assign out[2] = _U70_out;
assign out[1] = _U69_out;
assign out[0] = _U68_out;
endmodule

module array_delay_U54 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
wire [15:0] _U56_in;
wire _U56_clk;
wire [15:0] _U56_out;
wire [15:0] _U57_in;
wire _U57_clk;
wire [15:0] _U57_out;
wire [15:0] _U58_in;
wire _U58_clk;
wire [15:0] _U58_out;
wire [15:0] _U59_in;
wire _U59_clk;
wire [15:0] _U59_out;
assign _U55_in = in[0];
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign _U56_in = in[1];
assign _U56_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U56 (
    .in(_U56_in),
    .clk(_U56_clk),
    .out(_U56_out)
);
assign _U57_in = in[2];
assign _U57_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U57 (
    .in(_U57_in),
    .clk(_U57_clk),
    .out(_U57_out)
);
assign _U58_in = in[3];
assign _U58_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U58 (
    .in(_U58_in),
    .clk(_U58_clk),
    .out(_U58_out)
);
assign _U59_in = in[4];
assign _U59_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U59_in),
    .clk(_U59_clk),
    .out(_U59_out)
);
assign out[4] = _U59_out;
assign out[3] = _U58_out;
assign out[2] = _U57_out;
assign out[1] = _U56_out;
assign out[0] = _U55_out;
endmodule

module array_delay_U44 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U45_in;
wire _U45_clk;
wire [15:0] _U45_out;
wire [15:0] _U46_in;
wire _U46_clk;
wire [15:0] _U46_out;
wire [15:0] _U47_in;
wire _U47_clk;
wire [15:0] _U47_out;
wire [15:0] _U48_in;
wire _U48_clk;
wire [15:0] _U48_out;
wire [15:0] _U49_in;
wire _U49_clk;
wire [15:0] _U49_out;
assign _U45_in = in[0];
assign _U45_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U45 (
    .in(_U45_in),
    .clk(_U45_clk),
    .out(_U45_out)
);
assign _U46_in = in[1];
assign _U46_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(_U46_in),
    .clk(_U46_clk),
    .out(_U46_out)
);
assign _U47_in = in[2];
assign _U47_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U47 (
    .in(_U47_in),
    .clk(_U47_clk),
    .out(_U47_out)
);
assign _U48_in = in[3];
assign _U48_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U48 (
    .in(_U48_in),
    .clk(_U48_clk),
    .out(_U48_out)
);
assign _U49_in = in[4];
assign _U49_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U49_in),
    .clk(_U49_clk),
    .out(_U49_out)
);
assign out[4] = _U49_out;
assign out[3] = _U48_out;
assign out[2] = _U47_out;
assign out[1] = _U46_out;
assign out[0] = _U45_out;
endmodule

module array_delay_U31 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U32_in;
wire _U32_clk;
wire [15:0] _U32_out;
wire [15:0] _U33_in;
wire _U33_clk;
wire [15:0] _U33_out;
wire [15:0] _U34_in;
wire _U34_clk;
wire [15:0] _U34_out;
wire [15:0] _U35_in;
wire _U35_clk;
wire [15:0] _U35_out;
wire [15:0] _U36_in;
wire _U36_clk;
wire [15:0] _U36_out;
assign _U32_in = in[0];
assign _U32_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U32 (
    .in(_U32_in),
    .clk(_U32_clk),
    .out(_U32_out)
);
assign _U33_in = in[1];
assign _U33_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U33 (
    .in(_U33_in),
    .clk(_U33_clk),
    .out(_U33_out)
);
assign _U34_in = in[2];
assign _U34_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U34 (
    .in(_U34_in),
    .clk(_U34_clk),
    .out(_U34_out)
);
assign _U35_in = in[3];
assign _U35_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U35 (
    .in(_U35_in),
    .clk(_U35_clk),
    .out(_U35_out)
);
assign _U36_in = in[4];
assign _U36_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(_U36_in),
    .clk(_U36_clk),
    .out(_U36_out)
);
assign out[4] = _U36_out;
assign out[3] = _U35_out;
assign out[2] = _U34_out;
assign out[1] = _U33_out;
assign out[0] = _U32_out;
endmodule

module array_delay_U21 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U22_in;
wire _U22_clk;
wire [15:0] _U22_out;
wire [15:0] _U23_in;
wire _U23_clk;
wire [15:0] _U23_out;
wire [15:0] _U24_in;
wire _U24_clk;
wire [15:0] _U24_out;
wire [15:0] _U25_in;
wire _U25_clk;
wire [15:0] _U25_out;
wire [15:0] _U26_in;
wire _U26_clk;
wire [15:0] _U26_out;
assign _U22_in = in[0];
assign _U22_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U22 (
    .in(_U22_in),
    .clk(_U22_clk),
    .out(_U22_out)
);
assign _U23_in = in[1];
assign _U23_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U23 (
    .in(_U23_in),
    .clk(_U23_clk),
    .out(_U23_out)
);
assign _U24_in = in[2];
assign _U24_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U24 (
    .in(_U24_in),
    .clk(_U24_clk),
    .out(_U24_out)
);
assign _U25_in = in[3];
assign _U25_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U25 (
    .in(_U25_in),
    .clk(_U25_clk),
    .out(_U25_out)
);
assign _U26_in = in[4];
assign _U26_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U26 (
    .in(_U26_in),
    .clk(_U26_clk),
    .out(_U26_out)
);
assign out[4] = _U26_out;
assign out[3] = _U25_out;
assign out[2] = _U24_out;
assign out[1] = _U23_out;
assign out[0] = _U22_out;
endmodule

module array_delay_U105 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire _U108_clk;
wire [15:0] _U108_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
wire [15:0] _U110_in;
wire _U110_clk;
wire [15:0] _U110_out;
assign _U106_in = in[0];
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = in[1];
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = in[2];
assign _U108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U108_in),
    .clk(_U108_clk),
    .out(_U108_out)
);
assign _U109_in = in[3];
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign _U110_in = in[4];
assign _U110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U110_in),
    .clk(_U110_clk),
    .out(_U110_out)
);
assign out[4] = _U110_out;
assign out[3] = _U109_out;
assign out[2] = _U108_out;
assign out[1] = _U107_out;
assign out[0] = _U106_out;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U104_clk;
wire [15:0] arr__U104_in [4:0];
wire [15:0] arr__U104_out [4:0];
wire arr__U20_clk;
wire [15:0] arr__U20_in [4:0];
wire [15:0] arr__U20_out [4:0];
wire arr__U30_clk;
wire [15:0] arr__U30_in [4:0];
wire [15:0] arr__U30_out [4:0];
wire arr__U43_clk;
wire [15:0] arr__U43_in [4:0];
wire [15:0] arr__U43_out [4:0];
wire arr__U53_clk;
wire [15:0] arr__U53_in [4:0];
wire [15:0] arr__U53_out [4:0];
wire arr__U66_clk;
wire [15:0] arr__U66_in [3:0];
wire [15:0] arr__U66_out [3:0];
wire arr__U75_clk;
wire [15:0] arr__U75_in [3:0];
wire [15:0] arr__U75_out [3:0];
wire arr__U94_clk;
wire [15:0] arr__U94_in [4:0];
wire [15:0] arr__U94_out [4:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U102_clk;
wire delay_reg__U102_in;
wire delay_reg__U102_out;
wire delay_reg__U18_clk;
wire delay_reg__U18_in;
wire delay_reg__U18_out;
wire delay_reg__U28_clk;
wire delay_reg__U28_in;
wire delay_reg__U28_out;
wire delay_reg__U41_clk;
wire delay_reg__U41_in;
wire delay_reg__U41_out;
wire delay_reg__U51_clk;
wire delay_reg__U51_in;
wire delay_reg__U51_out;
wire delay_reg__U64_clk;
wire delay_reg__U64_in;
wire delay_reg__U64_out;
wire delay_reg__U73_clk;
wire delay_reg__U73_in;
wire delay_reg__U73_out;
wire delay_reg__U92_clk;
wire delay_reg__U92_in;
wire delay_reg__U92_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_rst_n;
wire op_hcompute_conv_stencil_1_port_controller_flush;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_rst_n;
wire op_hcompute_conv_stencil_2_port_controller_flush;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_rst_n;
wire op_hcompute_conv_stencil_3_port_controller_flush;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_rst_n;
wire op_hcompute_conv_stencil_4_port_controller_flush;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_rst_n;
wire op_hcompute_conv_stencil_5_port_controller_flush;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_rst_n;
wire op_hcompute_conv_stencil_port_controller_flush;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_rst_n;
wire op_hcompute_hw_output_stencil_port_controller_flush;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U104_clk = clk;
assign arr__U104_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U104_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U104_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U104_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U104_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U105 arr__U104 (
    .clk(arr__U104_clk),
    .in(arr__U104_in),
    .out(arr__U104_out)
);
assign arr__U20_clk = clk;
assign arr__U20_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U20_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U20_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U20_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U20_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U21 arr__U20 (
    .clk(arr__U20_clk),
    .in(arr__U20_in),
    .out(arr__U20_out)
);
assign arr__U30_clk = clk;
assign arr__U30_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U30_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U30_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U30_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U30_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U31 arr__U30 (
    .clk(arr__U30_clk),
    .in(arr__U30_in),
    .out(arr__U30_out)
);
assign arr__U43_clk = clk;
assign arr__U43_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U43_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U43_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U43_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U43_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U44 arr__U43 (
    .clk(arr__U43_clk),
    .in(arr__U43_in),
    .out(arr__U43_out)
);
assign arr__U53_clk = clk;
assign arr__U53_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U53_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U53_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U53_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U53_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U54 arr__U53 (
    .clk(arr__U53_clk),
    .in(arr__U53_in),
    .out(arr__U53_out)
);
assign arr__U66_clk = clk;
assign arr__U66_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U66_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U66_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U66_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U67 arr__U66 (
    .clk(arr__U66_clk),
    .in(arr__U66_in),
    .out(arr__U66_out)
);
assign arr__U75_clk = clk;
assign arr__U75_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U75_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U75_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U75_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U76 arr__U75 (
    .clk(arr__U75_clk),
    .in(arr__U75_in),
    .out(arr__U75_out)
);
assign arr__U94_clk = clk;
assign arr__U94_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U94_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U94_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U94_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U94_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U95 arr__U94 (
    .clk(arr__U94_clk),
    .in(arr__U94_in),
    .out(arr__U94_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U102_clk = clk;
assign delay_reg__U102_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U102 (
    .clk(delay_reg__U102_clk),
    .in(delay_reg__U102_in),
    .out(delay_reg__U102_out)
);
assign delay_reg__U18_clk = clk;
assign delay_reg__U18_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U18 (
    .clk(delay_reg__U18_clk),
    .in(delay_reg__U18_in),
    .out(delay_reg__U18_out)
);
assign delay_reg__U28_clk = clk;
assign delay_reg__U28_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U28 (
    .clk(delay_reg__U28_clk),
    .in(delay_reg__U28_in),
    .out(delay_reg__U28_out)
);
assign delay_reg__U41_clk = clk;
assign delay_reg__U41_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U41 (
    .clk(delay_reg__U41_clk),
    .in(delay_reg__U41_in),
    .out(delay_reg__U41_out)
);
assign delay_reg__U51_clk = clk;
assign delay_reg__U51_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U51 (
    .clk(delay_reg__U51_clk),
    .in(delay_reg__U51_in),
    .out(delay_reg__U51_out)
);
assign delay_reg__U64_clk = clk;
assign delay_reg__U64_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U64 (
    .clk(delay_reg__U64_clk),
    .in(delay_reg__U64_in),
    .out(delay_reg__U64_out)
);
assign delay_reg__U73_clk = clk;
assign delay_reg__U73_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U73 (
    .clk(delay_reg__U73_clk),
    .in(delay_reg__U73_in),
    .out(delay_reg__U73_out)
);
assign delay_reg__U92_clk = clk;
assign delay_reg__U92_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U92 (
    .clk(delay_reg__U92_clk),
    .in(delay_reg__U92_in),
    .out(delay_reg__U92_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U3 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U4 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
assign op_hcompute_conv_stencil_1_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_1_port_controller_flush = flush;
affine_controller__U0 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_1_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_1_port_controller_flush),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U1 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U2 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U5 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U6 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U10 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U11 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
assign op_hcompute_conv_stencil_2_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_2_port_controller_flush = flush;
affine_controller__U7 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_2_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_2_port_controller_flush),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U8 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U9 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U12 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U13 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U92_out;
op_hcompute_conv_stencil_3_exe_start_pt__U91 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U94_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U94_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U94_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U94_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U94_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U93 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
assign op_hcompute_conv_stencil_3_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_3_port_controller_flush = flush;
affine_controller__U88 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_3_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_3_port_controller_flush),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U89 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U90 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U102_out;
op_hcompute_conv_stencil_3_write_start_pt__U101 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U104_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U104_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U104_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U104_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U104_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U103 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U18_out;
op_hcompute_conv_stencil_4_exe_start_pt__U17 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U20_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U20_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U20_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U20_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U20_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U19 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
assign op_hcompute_conv_stencil_4_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_4_port_controller_flush = flush;
affine_controller__U14 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_4_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_4_port_controller_flush),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U15 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U16 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U28_out;
op_hcompute_conv_stencil_4_write_start_pt__U27 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U30_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U30_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U30_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U30_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U30_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U29 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U41_out;
op_hcompute_conv_stencil_5_exe_start_pt__U40 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U43_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U43_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U43_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U43_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U43_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U42 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
assign op_hcompute_conv_stencil_5_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_5_port_controller_flush = flush;
affine_controller__U37 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_5_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_5_port_controller_flush),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U38 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U39 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U51_out;
op_hcompute_conv_stencil_5_write_start_pt__U50 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U53_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U53_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U53_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U53_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U53_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U52 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U121 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U122 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
assign op_hcompute_conv_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_port_controller_flush = flush;
affine_controller__U118 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_port_controller_flush),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U119 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U120 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U123 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U124 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U84 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U85 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U81 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U82 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U83 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U86 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U87 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U114 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U115 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U111 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U112 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U113 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U116 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U117 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U64_out;
op_hcompute_hw_output_stencil_exe_start_pt__U63 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U66_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U66_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U66_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U66_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U65 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
assign op_hcompute_hw_output_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_output_stencil_port_controller_flush = flush;
affine_controller__U60 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_output_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_output_stencil_port_controller_flush),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U61 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U62 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U73_out;
op_hcompute_hw_output_stencil_write_start_pt__U72 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U75_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U75_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U75_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U75_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U74 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

