// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
// Module `affine_controller__U81` defined externally
// Module `affine_controller__U74` defined externally
// Module `affine_controller__U51` defined externally
// Module `affine_controller__U44` defined externally
// Module `affine_controller__U37` defined externally
// Module `affine_controller__U30` defined externally
// Module `affine_controller__U23` defined externally
// Module `affine_controller__U102` defined externally
// Module `affine_controller__U0` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U93 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U95 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U82 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U83 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U84 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U86 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U42 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U43 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U38 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U39 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U41 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U79 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U80 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U75 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U76 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U77 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U78 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U49 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U50 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U45 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U46 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U47 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U48 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U13 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U15 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U1 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U2 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U3 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U5 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U64 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U66 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U52 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U53 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U54 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U56 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U115 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U117 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U103 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U104 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U105 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U107 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U35 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U36 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U31 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U32 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U33 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U34 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U28 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U29 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U24 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U25 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U26 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U27 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module hcompute_hw_output_stencil (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
assign out_hw_output_stencil = in0_conv_stencil[0];
endmodule

module hcompute_hw_kernel_global_wrapper_stencil (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
assign out_hw_kernel_global_wrapper_stencil = in0_hw_kernel_stencil[0];
endmodule

module hcompute_hw_input_global_wrapper_stencil (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
assign out_hw_input_global_wrapper_stencil = in0_hw_input_stencil[0];
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module hcompute_conv_stencil_2 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_1 (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil (
    output [15:0] out_conv_stencil
);
assign out_conv_stencil = 16'h0000;
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_5 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_4 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module hcompute_conv_stencil_3 (
    output [15:0] out_conv_stencil,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0]
);
assign out_conv_stencil = 16'((16'(in2_hw_kernel_global_wrapper_stencil[0] * in1_hw_input_global_wrapper_stencil[0])) + (16'(in0_conv_stencil[0] + (16'((16'(in2_hw_kernel_global_wrapper_stencil[1] * in1_hw_input_global_wrapper_stencil[1])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[2] * in1_hw_input_global_wrapper_stencil[2])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[3] * in1_hw_input_global_wrapper_stencil[3])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[4] * in1_hw_input_global_wrapper_stencil[4])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[5] * in1_hw_input_global_wrapper_stencil[5])) + (16'((16'(in2_hw_kernel_global_wrapper_stencil[6] * in1_hw_input_global_wrapper_stencil[6])) + (16'(in2_hw_kernel_global_wrapper_stencil[7] * in1_hw_input_global_wrapper_stencil[7])))))))))))))))));
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3 inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U97 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U100_in = in[2];
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = in[3];
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U98_in = in[0];
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = in[1];
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
assign out[3] = _U101_out;
assign out[2] = _U100_out;
assign out[1] = _U99_out;
assign out[0] = _U98_out;
endmodule

module array_delay_U88 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U89_in;
wire _U89_clk;
wire [15:0] _U89_out;
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
assign _U89_in = in[0];
assign _U89_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U89 (
    .in(_U89_in),
    .clk(_U89_clk),
    .out(_U89_out)
);
assign _U90_in = in[1];
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = in[2];
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = in[3];
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign out[3] = _U92_out;
assign out[2] = _U91_out;
assign out[1] = _U90_out;
assign out[0] = _U89_out;
endmodule

module array_delay_U7 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U10_in;
wire _U10_clk;
wire [15:0] _U10_out;
wire [15:0] _U11_in;
wire _U11_clk;
wire [15:0] _U11_out;
wire [15:0] _U12_in;
wire _U12_clk;
wire [15:0] _U12_out;
wire [15:0] _U8_in;
wire _U8_clk;
wire [15:0] _U8_out;
wire [15:0] _U9_in;
wire _U9_clk;
wire [15:0] _U9_out;
assign _U10_in = in[2];
assign _U10_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U10 (
    .in(_U10_in),
    .clk(_U10_clk),
    .out(_U10_out)
);
assign _U11_in = in[3];
assign _U11_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U11 (
    .in(_U11_in),
    .clk(_U11_clk),
    .out(_U11_out)
);
assign _U12_in = in[4];
assign _U12_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U12 (
    .in(_U12_in),
    .clk(_U12_clk),
    .out(_U12_out)
);
assign _U8_in = in[0];
assign _U8_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U8 (
    .in(_U8_in),
    .clk(_U8_clk),
    .out(_U8_out)
);
assign _U9_in = in[1];
assign _U9_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U9 (
    .in(_U9_in),
    .clk(_U9_clk),
    .out(_U9_out)
);
assign out[4] = _U12_out;
assign out[3] = _U11_out;
assign out[2] = _U10_out;
assign out[1] = _U9_out;
assign out[0] = _U8_out;
endmodule

module array_delay_U68 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U69_in;
wire _U69_clk;
wire [15:0] _U69_out;
wire [15:0] _U70_in;
wire _U70_clk;
wire [15:0] _U70_out;
wire [15:0] _U71_in;
wire _U71_clk;
wire [15:0] _U71_out;
wire [15:0] _U72_in;
wire _U72_clk;
wire [15:0] _U72_out;
wire [15:0] _U73_in;
wire _U73_clk;
wire [15:0] _U73_out;
assign _U69_in = in[0];
assign _U69_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(_U69_in),
    .clk(_U69_clk),
    .out(_U69_out)
);
assign _U70_in = in[1];
assign _U70_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U70 (
    .in(_U70_in),
    .clk(_U70_clk),
    .out(_U70_out)
);
assign _U71_in = in[2];
assign _U71_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U71 (
    .in(_U71_in),
    .clk(_U71_clk),
    .out(_U71_out)
);
assign _U72_in = in[3];
assign _U72_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U72 (
    .in(_U72_in),
    .clk(_U72_clk),
    .out(_U72_out)
);
assign _U73_in = in[4];
assign _U73_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U73 (
    .in(_U73_in),
    .clk(_U73_clk),
    .out(_U73_out)
);
assign out[4] = _U73_out;
assign out[3] = _U72_out;
assign out[2] = _U71_out;
assign out[1] = _U70_out;
assign out[0] = _U69_out;
endmodule

module array_delay_U58 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U59_in;
wire _U59_clk;
wire [15:0] _U59_out;
wire [15:0] _U60_in;
wire _U60_clk;
wire [15:0] _U60_out;
wire [15:0] _U61_in;
wire _U61_clk;
wire [15:0] _U61_out;
wire [15:0] _U62_in;
wire _U62_clk;
wire [15:0] _U62_out;
wire [15:0] _U63_in;
wire _U63_clk;
wire [15:0] _U63_out;
assign _U59_in = in[0];
assign _U59_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U59_in),
    .clk(_U59_clk),
    .out(_U59_out)
);
assign _U60_in = in[1];
assign _U60_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U60 (
    .in(_U60_in),
    .clk(_U60_clk),
    .out(_U60_out)
);
assign _U61_in = in[2];
assign _U61_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U61 (
    .in(_U61_in),
    .clk(_U61_clk),
    .out(_U61_out)
);
assign _U62_in = in[3];
assign _U62_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U62 (
    .in(_U62_in),
    .clk(_U62_clk),
    .out(_U62_out)
);
assign _U63_in = in[4];
assign _U63_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U63 (
    .in(_U63_in),
    .clk(_U63_clk),
    .out(_U63_out)
);
assign out[4] = _U63_out;
assign out[3] = _U62_out;
assign out[2] = _U61_out;
assign out[1] = _U60_out;
assign out[0] = _U59_out;
endmodule

module array_delay_U17 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U18_in;
wire _U18_clk;
wire [15:0] _U18_out;
wire [15:0] _U19_in;
wire _U19_clk;
wire [15:0] _U19_out;
wire [15:0] _U20_in;
wire _U20_clk;
wire [15:0] _U20_out;
wire [15:0] _U21_in;
wire _U21_clk;
wire [15:0] _U21_out;
wire [15:0] _U22_in;
wire _U22_clk;
wire [15:0] _U22_out;
assign _U18_in = in[0];
assign _U18_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U18 (
    .in(_U18_in),
    .clk(_U18_clk),
    .out(_U18_out)
);
assign _U19_in = in[1];
assign _U19_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U19 (
    .in(_U19_in),
    .clk(_U19_clk),
    .out(_U19_out)
);
assign _U20_in = in[2];
assign _U20_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U20 (
    .in(_U20_in),
    .clk(_U20_clk),
    .out(_U20_out)
);
assign _U21_in = in[3];
assign _U21_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U21 (
    .in(_U21_in),
    .clk(_U21_clk),
    .out(_U21_out)
);
assign _U22_in = in[4];
assign _U22_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U22 (
    .in(_U22_in),
    .clk(_U22_clk),
    .out(_U22_out)
);
assign out[4] = _U22_out;
assign out[3] = _U21_out;
assign out[2] = _U20_out;
assign out[1] = _U19_out;
assign out[0] = _U18_out;
endmodule

module array_delay_U119 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U120_in;
wire _U120_clk;
wire [15:0] _U120_out;
wire [15:0] _U121_in;
wire _U121_clk;
wire [15:0] _U121_out;
wire [15:0] _U122_in;
wire _U122_clk;
wire [15:0] _U122_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
assign _U120_in = in[0];
assign _U120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(_U120_in),
    .clk(_U120_clk),
    .out(_U120_out)
);
assign _U121_in = in[1];
assign _U121_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U121 (
    .in(_U121_in),
    .clk(_U121_clk),
    .out(_U121_out)
);
assign _U122_in = in[2];
assign _U122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U122 (
    .in(_U122_in),
    .clk(_U122_clk),
    .out(_U122_out)
);
assign _U123_in = in[3];
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = in[4];
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign out[4] = _U124_out;
assign out[3] = _U123_out;
assign out[2] = _U122_out;
assign out[1] = _U121_out;
assign out[0] = _U120_out;
endmodule

module array_delay_U109 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U110_in;
wire _U110_clk;
wire [15:0] _U110_out;
wire [15:0] _U111_in;
wire _U111_clk;
wire [15:0] _U111_out;
wire [15:0] _U112_in;
wire _U112_clk;
wire [15:0] _U112_out;
wire [15:0] _U113_in;
wire _U113_clk;
wire [15:0] _U113_out;
wire [15:0] _U114_in;
wire _U114_clk;
wire [15:0] _U114_out;
assign _U110_in = in[0];
assign _U110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U110_in),
    .clk(_U110_clk),
    .out(_U110_out)
);
assign _U111_in = in[1];
assign _U111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U111 (
    .in(_U111_in),
    .clk(_U111_clk),
    .out(_U111_out)
);
assign _U112_in = in[2];
assign _U112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U112_in),
    .clk(_U112_clk),
    .out(_U112_out)
);
assign _U113_in = in[3];
assign _U113_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U113 (
    .in(_U113_in),
    .clk(_U113_clk),
    .out(_U113_out)
);
assign _U114_in = in[4];
assign _U114_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U114 (
    .in(_U114_in),
    .clk(_U114_clk),
    .out(_U114_out)
);
assign out[4] = _U114_out;
assign out[3] = _U113_out;
assign out[2] = _U112_out;
assign out[1] = _U111_out;
assign out[0] = _U110_out;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U108_clk;
wire [15:0] arr__U108_in [4:0];
wire [15:0] arr__U108_out [4:0];
wire arr__U118_clk;
wire [15:0] arr__U118_in [4:0];
wire [15:0] arr__U118_out [4:0];
wire arr__U16_clk;
wire [15:0] arr__U16_in [4:0];
wire [15:0] arr__U16_out [4:0];
wire arr__U57_clk;
wire [15:0] arr__U57_in [4:0];
wire [15:0] arr__U57_out [4:0];
wire arr__U6_clk;
wire [15:0] arr__U6_in [4:0];
wire [15:0] arr__U6_out [4:0];
wire arr__U67_clk;
wire [15:0] arr__U67_in [4:0];
wire [15:0] arr__U67_out [4:0];
wire arr__U87_clk;
wire [15:0] arr__U87_in [3:0];
wire [15:0] arr__U87_out [3:0];
wire arr__U96_clk;
wire [15:0] arr__U96_in [3:0];
wire [15:0] arr__U96_out [3:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U106_clk;
wire delay_reg__U106_in;
wire delay_reg__U106_out;
wire delay_reg__U116_clk;
wire delay_reg__U116_in;
wire delay_reg__U116_out;
wire delay_reg__U14_clk;
wire delay_reg__U14_in;
wire delay_reg__U14_out;
wire delay_reg__U4_clk;
wire delay_reg__U4_in;
wire delay_reg__U4_out;
wire delay_reg__U55_clk;
wire delay_reg__U55_in;
wire delay_reg__U55_out;
wire delay_reg__U65_clk;
wire delay_reg__U65_in;
wire delay_reg__U65_out;
wire delay_reg__U85_clk;
wire delay_reg__U85_in;
wire delay_reg__U85_out;
wire delay_reg__U94_clk;
wire delay_reg__U94_in;
wire delay_reg__U94_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_rst_n;
wire op_hcompute_conv_stencil_1_port_controller_flush;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_rst_n;
wire op_hcompute_conv_stencil_2_port_controller_flush;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_rst_n;
wire op_hcompute_conv_stencil_3_port_controller_flush;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_rst_n;
wire op_hcompute_conv_stencil_4_port_controller_flush;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_rst_n;
wire op_hcompute_conv_stencil_5_port_controller_flush;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_rst_n;
wire op_hcompute_conv_stencil_port_controller_flush;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_rst_n;
wire op_hcompute_hw_output_stencil_port_controller_flush;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U108_clk = clk;
assign arr__U108_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U108_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U108_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U108_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U108_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U109 arr__U108 (
    .clk(arr__U108_clk),
    .in(arr__U108_in),
    .out(arr__U108_out)
);
assign arr__U118_clk = clk;
assign arr__U118_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U118_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U118_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U118_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U118_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U119 arr__U118 (
    .clk(arr__U118_clk),
    .in(arr__U118_in),
    .out(arr__U118_out)
);
assign arr__U16_clk = clk;
assign arr__U16_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U16_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U16_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U16_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U16_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U17 arr__U16 (
    .clk(arr__U16_clk),
    .in(arr__U16_in),
    .out(arr__U16_out)
);
assign arr__U57_clk = clk;
assign arr__U57_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U57_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U57_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U57_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U57_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U58 arr__U57 (
    .clk(arr__U57_clk),
    .in(arr__U57_in),
    .out(arr__U57_out)
);
assign arr__U6_clk = clk;
assign arr__U6_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U6_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U6_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U6_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U6_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U7 arr__U6 (
    .clk(arr__U6_clk),
    .in(arr__U6_in),
    .out(arr__U6_out)
);
assign arr__U67_clk = clk;
assign arr__U67_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U67_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U67_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U67_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U67_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U68 arr__U67 (
    .clk(arr__U67_clk),
    .in(arr__U67_in),
    .out(arr__U67_out)
);
assign arr__U87_clk = clk;
assign arr__U87_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U87_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U87_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U87_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U88 arr__U87 (
    .clk(arr__U87_clk),
    .in(arr__U87_in),
    .out(arr__U87_out)
);
assign arr__U96_clk = clk;
assign arr__U96_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U96_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U96_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U96_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U97 arr__U96 (
    .clk(arr__U96_clk),
    .in(arr__U96_in),
    .out(arr__U96_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U106_clk = clk;
assign delay_reg__U106_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U106 (
    .clk(delay_reg__U106_clk),
    .in(delay_reg__U106_in),
    .out(delay_reg__U106_out)
);
assign delay_reg__U116_clk = clk;
assign delay_reg__U116_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U116 (
    .clk(delay_reg__U116_clk),
    .in(delay_reg__U116_in),
    .out(delay_reg__U116_out)
);
assign delay_reg__U14_clk = clk;
assign delay_reg__U14_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U14 (
    .clk(delay_reg__U14_clk),
    .in(delay_reg__U14_in),
    .out(delay_reg__U14_out)
);
assign delay_reg__U4_clk = clk;
assign delay_reg__U4_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U4 (
    .clk(delay_reg__U4_clk),
    .in(delay_reg__U4_in),
    .out(delay_reg__U4_out)
);
assign delay_reg__U55_clk = clk;
assign delay_reg__U55_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U55 (
    .clk(delay_reg__U55_clk),
    .in(delay_reg__U55_in),
    .out(delay_reg__U55_out)
);
assign delay_reg__U65_clk = clk;
assign delay_reg__U65_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U65 (
    .clk(delay_reg__U65_clk),
    .in(delay_reg__U65_in),
    .out(delay_reg__U65_out)
);
assign delay_reg__U85_clk = clk;
assign delay_reg__U85_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U85 (
    .clk(delay_reg__U85_clk),
    .in(delay_reg__U85_in),
    .out(delay_reg__U85_out)
);
assign delay_reg__U94_clk = clk;
assign delay_reg__U94_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U94 (
    .clk(delay_reg__U94_clk),
    .in(delay_reg__U94_in),
    .out(delay_reg__U94_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U26 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U27 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
assign op_hcompute_conv_stencil_1_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_1_port_controller_flush = flush;
affine_controller__U23 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_1_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_1_port_controller_flush),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U24 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U25 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U28 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U29 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U33 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U34 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
assign op_hcompute_conv_stencil_2_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_2_port_controller_flush = flush;
affine_controller__U30 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_2_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_2_port_controller_flush),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U31 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U32 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U35 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U36 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U106_out;
op_hcompute_conv_stencil_3_exe_start_pt__U105 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U108_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U108_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U108_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U108_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U108_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U107 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
assign op_hcompute_conv_stencil_3_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_3_port_controller_flush = flush;
affine_controller__U102 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_3_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_3_port_controller_flush),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U103 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U104 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U116_out;
op_hcompute_conv_stencil_3_write_start_pt__U115 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U118_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U118_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U118_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U118_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U118_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U117 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U55_out;
op_hcompute_conv_stencil_4_exe_start_pt__U54 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U57_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U57_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U57_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U57_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U57_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U56 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
assign op_hcompute_conv_stencil_4_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_4_port_controller_flush = flush;
affine_controller__U51 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_4_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_4_port_controller_flush),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U52 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U53 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U65_out;
op_hcompute_conv_stencil_4_write_start_pt__U64 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U67_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U67_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U67_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U67_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U67_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U66 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U4_out;
op_hcompute_conv_stencil_5_exe_start_pt__U3 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U6_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U6_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U6_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U6_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U6_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U5 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
assign op_hcompute_conv_stencil_5_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_5_port_controller_flush = flush;
affine_controller__U0 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_5_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_5_port_controller_flush),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U1 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U2 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U14_out;
op_hcompute_conv_stencil_5_write_start_pt__U13 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U16_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U16_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U16_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U16_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U16_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U15 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U47 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U48 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
assign op_hcompute_conv_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_port_controller_flush = flush;
affine_controller__U44 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_port_controller_flush),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U45 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U46 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U49 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U50 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U77 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U78 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U74 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U75 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U76 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U79 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U80 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U40 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U41 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U37 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U38 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U39 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U42 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U43 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U85_out;
op_hcompute_hw_output_stencil_exe_start_pt__U84 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U87_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U87_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U87_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U87_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U86 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
assign op_hcompute_hw_output_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_output_stencil_port_controller_flush = flush;
affine_controller__U81 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_output_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_output_stencil_port_controller_flush),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U82 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U83 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U94_out;
op_hcompute_hw_output_stencil_write_start_pt__U93 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U96_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U96_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U96_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U96_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U95 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

