// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
// Module `affine_controller__U7` defined externally
// Module `affine_controller__U63` defined externally
// Module `affine_controller__U56` defined externally
// Module `affine_controller__U388` defined externally
// Module `affine_controller__U381` defined externally
// Module `affine_controller__U222` defined externally
// Module `affine_controller__U21` defined externally
// Module `affine_controller__U14` defined externally
// Module `affine_controller__U0` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U43 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U22 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U23 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U24 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U27 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U61 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U62 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U57 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U58 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U59 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U60 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U5 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U6 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U1 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U2 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U3 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U4 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U19 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U20 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U15 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U16 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U17 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U18 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U243 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U261 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U223 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U224 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U225 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U228 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U84 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U102 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U64 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U65 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U66 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U69 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U409 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U427 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U389 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U390 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U391 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U394 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U386 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U387 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U382 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U383 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U384 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U385 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U12 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U13 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U8 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U9 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U10 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U11 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U78 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U79_in;
wire _U79_clk;
wire [15:0] _U79_out;
wire [15:0] _U80_in;
wire _U80_clk;
wire [15:0] _U80_out;
wire [15:0] _U81_in;
wire _U81_clk;
wire [15:0] _U81_out;
wire [15:0] _U82_in;
wire _U82_clk;
wire [15:0] _U82_out;
wire [15:0] _U83_in;
wire _U83_clk;
wire [15:0] _U83_out;
assign _U79_in = in[0];
assign _U79_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(_U79_in),
    .clk(_U79_clk),
    .out(_U79_out)
);
assign _U80_in = in[1];
assign _U80_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(_U80_in),
    .clk(_U80_clk),
    .out(_U80_out)
);
assign _U81_in = in[2];
assign _U81_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U81 (
    .in(_U81_in),
    .clk(_U81_clk),
    .out(_U81_out)
);
assign _U82_in = in[3];
assign _U82_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U82 (
    .in(_U82_in),
    .clk(_U82_clk),
    .out(_U82_out)
);
assign _U83_in = in[4];
assign _U83_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U83 (
    .in(_U83_in),
    .clk(_U83_clk),
    .out(_U83_out)
);
assign out[4] = _U83_out;
assign out[3] = _U82_out;
assign out[2] = _U81_out;
assign out[1] = _U80_out;
assign out[0] = _U79_out;
endmodule

module array_delay_U71 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U72_in;
wire _U72_clk;
wire [15:0] _U72_out;
wire [15:0] _U73_in;
wire _U73_clk;
wire [15:0] _U73_out;
wire [15:0] _U74_in;
wire _U74_clk;
wire [15:0] _U74_out;
wire [15:0] _U75_in;
wire _U75_clk;
wire [15:0] _U75_out;
wire [15:0] _U76_in;
wire _U76_clk;
wire [15:0] _U76_out;
assign _U72_in = in[0];
assign _U72_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U72 (
    .in(_U72_in),
    .clk(_U72_clk),
    .out(_U72_out)
);
assign _U73_in = in[1];
assign _U73_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U73 (
    .in(_U73_in),
    .clk(_U73_clk),
    .out(_U73_out)
);
assign _U74_in = in[2];
assign _U74_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U74 (
    .in(_U74_in),
    .clk(_U74_clk),
    .out(_U74_out)
);
assign _U75_in = in[3];
assign _U75_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U75 (
    .in(_U75_in),
    .clk(_U75_clk),
    .out(_U75_out)
);
assign _U76_in = in[4];
assign _U76_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U76 (
    .in(_U76_in),
    .clk(_U76_clk),
    .out(_U76_out)
);
assign out[4] = _U76_out;
assign out[3] = _U75_out;
assign out[2] = _U74_out;
assign out[1] = _U73_out;
assign out[0] = _U72_out;
endmodule

module array_delay_U541 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
wire [15:0] _U543_in;
wire _U543_clk;
wire [15:0] _U543_out;
wire [15:0] _U544_in;
wire _U544_clk;
wire [15:0] _U544_out;
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
assign _U542_in = in[0];
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign _U543_in = in[1];
assign _U543_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U543 (
    .in(_U543_in),
    .clk(_U543_clk),
    .out(_U543_out)
);
assign _U544_in = in[2];
assign _U544_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U544 (
    .in(_U544_in),
    .clk(_U544_clk),
    .out(_U544_out)
);
assign _U545_in = in[3];
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = in[4];
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign out[4] = _U546_out;
assign out[3] = _U545_out;
assign out[2] = _U544_out;
assign out[1] = _U543_out;
assign out[0] = _U542_out;
endmodule

module array_delay_U534 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U535_in;
wire _U535_clk;
wire [15:0] _U535_out;
wire [15:0] _U536_in;
wire _U536_clk;
wire [15:0] _U536_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire _U539_clk;
wire [15:0] _U539_out;
assign _U535_in = in[0];
assign _U535_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(_U535_in),
    .clk(_U535_clk),
    .out(_U535_out)
);
assign _U536_in = in[1];
assign _U536_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U536_in),
    .clk(_U536_clk),
    .out(_U536_out)
);
assign _U537_in = in[2];
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign _U538_in = in[3];
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = in[4];
assign _U539_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U539_in),
    .clk(_U539_clk),
    .out(_U539_out)
);
assign out[4] = _U539_out;
assign out[3] = _U538_out;
assign out[2] = _U537_out;
assign out[1] = _U536_out;
assign out[0] = _U535_out;
endmodule

module array_delay_U527 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U528_in;
wire _U528_clk;
wire [15:0] _U528_out;
wire [15:0] _U529_in;
wire _U529_clk;
wire [15:0] _U529_out;
wire [15:0] _U530_in;
wire _U530_clk;
wire [15:0] _U530_out;
wire [15:0] _U531_in;
wire _U531_clk;
wire [15:0] _U531_out;
wire [15:0] _U532_in;
wire _U532_clk;
wire [15:0] _U532_out;
assign _U528_in = in[0];
assign _U528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(_U528_in),
    .clk(_U528_clk),
    .out(_U528_out)
);
assign _U529_in = in[1];
assign _U529_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U529 (
    .in(_U529_in),
    .clk(_U529_clk),
    .out(_U529_out)
);
assign _U530_in = in[2];
assign _U530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U530 (
    .in(_U530_in),
    .clk(_U530_clk),
    .out(_U530_out)
);
assign _U531_in = in[3];
assign _U531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(_U531_in),
    .clk(_U531_clk),
    .out(_U531_out)
);
assign _U532_in = in[4];
assign _U532_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U532 (
    .in(_U532_in),
    .clk(_U532_clk),
    .out(_U532_out)
);
assign out[4] = _U532_out;
assign out[3] = _U531_out;
assign out[2] = _U530_out;
assign out[1] = _U529_out;
assign out[0] = _U528_out;
endmodule

module array_delay_U520 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U521_in;
wire _U521_clk;
wire [15:0] _U521_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
wire [15:0] _U524_in;
wire _U524_clk;
wire [15:0] _U524_out;
wire [15:0] _U525_in;
wire _U525_clk;
wire [15:0] _U525_out;
assign _U521_in = in[0];
assign _U521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U521_in),
    .clk(_U521_clk),
    .out(_U521_out)
);
assign _U522_in = in[1];
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = in[2];
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign _U524_in = in[3];
assign _U524_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U524 (
    .in(_U524_in),
    .clk(_U524_clk),
    .out(_U524_out)
);
assign _U525_in = in[4];
assign _U525_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U525 (
    .in(_U525_in),
    .clk(_U525_clk),
    .out(_U525_out)
);
assign out[4] = _U525_out;
assign out[3] = _U524_out;
assign out[2] = _U523_out;
assign out[1] = _U522_out;
assign out[0] = _U521_out;
endmodule

module array_delay_U513 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
wire [15:0] _U517_in;
wire _U517_clk;
wire [15:0] _U517_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
assign _U514_in = in[0];
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = in[1];
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = in[2];
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign _U517_in = in[3];
assign _U517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(_U517_in),
    .clk(_U517_clk),
    .out(_U517_out)
);
assign _U518_in = in[4];
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign out[4] = _U518_out;
assign out[3] = _U517_out;
assign out[2] = _U516_out;
assign out[1] = _U515_out;
assign out[0] = _U514_out;
endmodule

module array_delay_U51 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U52_in;
wire _U52_clk;
wire [15:0] _U52_out;
wire [15:0] _U53_in;
wire _U53_clk;
wire [15:0] _U53_out;
wire [15:0] _U54_in;
wire _U54_clk;
wire [15:0] _U54_out;
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
assign _U52_in = in[0];
assign _U52_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U52 (
    .in(_U52_in),
    .clk(_U52_clk),
    .out(_U52_out)
);
assign _U53_in = in[1];
assign _U53_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U53 (
    .in(_U53_in),
    .clk(_U53_clk),
    .out(_U53_out)
);
assign _U54_in = in[2];
assign _U54_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U54 (
    .in(_U54_in),
    .clk(_U54_clk),
    .out(_U54_out)
);
assign _U55_in = in[3];
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign out[3] = _U55_out;
assign out[2] = _U54_out;
assign out[1] = _U53_out;
assign out[0] = _U52_out;
endmodule

module array_delay_U506 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U507_in;
wire _U507_clk;
wire [15:0] _U507_out;
wire [15:0] _U508_in;
wire _U508_clk;
wire [15:0] _U508_out;
wire [15:0] _U509_in;
wire _U509_clk;
wire [15:0] _U509_out;
wire [15:0] _U510_in;
wire _U510_clk;
wire [15:0] _U510_out;
wire [15:0] _U511_in;
wire _U511_clk;
wire [15:0] _U511_out;
assign _U507_in = in[0];
assign _U507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U507 (
    .in(_U507_in),
    .clk(_U507_clk),
    .out(_U507_out)
);
assign _U508_in = in[1];
assign _U508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U508 (
    .in(_U508_in),
    .clk(_U508_clk),
    .out(_U508_out)
);
assign _U509_in = in[2];
assign _U509_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U509 (
    .in(_U509_in),
    .clk(_U509_clk),
    .out(_U509_out)
);
assign _U510_in = in[3];
assign _U510_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U510 (
    .in(_U510_in),
    .clk(_U510_clk),
    .out(_U510_out)
);
assign _U511_in = in[4];
assign _U511_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(_U511_in),
    .clk(_U511_clk),
    .out(_U511_out)
);
assign out[4] = _U511_out;
assign out[3] = _U510_out;
assign out[2] = _U509_out;
assign out[1] = _U508_out;
assign out[0] = _U507_out;
endmodule

module array_delay_U499 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire _U502_clk;
wire [15:0] _U502_out;
wire [15:0] _U503_in;
wire _U503_clk;
wire [15:0] _U503_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
assign _U500_in = in[0];
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign _U501_in = in[1];
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = in[2];
assign _U502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U502_in),
    .clk(_U502_clk),
    .out(_U502_out)
);
assign _U503_in = in[3];
assign _U503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(_U503_in),
    .clk(_U503_clk),
    .out(_U503_out)
);
assign _U504_in = in[4];
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign out[4] = _U504_out;
assign out[3] = _U503_out;
assign out[2] = _U502_out;
assign out[1] = _U501_out;
assign out[0] = _U500_out;
endmodule

module array_delay_U492 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U493_in;
wire _U493_clk;
wire [15:0] _U493_out;
wire [15:0] _U494_in;
wire _U494_clk;
wire [15:0] _U494_out;
wire [15:0] _U495_in;
wire _U495_clk;
wire [15:0] _U495_out;
wire [15:0] _U496_in;
wire _U496_clk;
wire [15:0] _U496_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
assign _U493_in = in[0];
assign _U493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U493 (
    .in(_U493_in),
    .clk(_U493_clk),
    .out(_U493_out)
);
assign _U494_in = in[1];
assign _U494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U494 (
    .in(_U494_in),
    .clk(_U494_clk),
    .out(_U494_out)
);
assign _U495_in = in[2];
assign _U495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U495 (
    .in(_U495_in),
    .clk(_U495_clk),
    .out(_U495_out)
);
assign _U496_in = in[3];
assign _U496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(_U496_in),
    .clk(_U496_clk),
    .out(_U496_out)
);
assign _U497_in = in[4];
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign out[4] = _U497_out;
assign out[3] = _U496_out;
assign out[2] = _U495_out;
assign out[1] = _U494_out;
assign out[0] = _U493_out;
endmodule

module array_delay_U485 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire _U487_clk;
wire [15:0] _U487_out;
wire [15:0] _U488_in;
wire _U488_clk;
wire [15:0] _U488_out;
wire [15:0] _U489_in;
wire _U489_clk;
wire [15:0] _U489_out;
wire [15:0] _U490_in;
wire _U490_clk;
wire [15:0] _U490_out;
assign _U486_in = in[0];
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = in[1];
assign _U487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U487 (
    .in(_U487_in),
    .clk(_U487_clk),
    .out(_U487_out)
);
assign _U488_in = in[2];
assign _U488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U488 (
    .in(_U488_in),
    .clk(_U488_clk),
    .out(_U488_out)
);
assign _U489_in = in[3];
assign _U489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U489_in),
    .clk(_U489_clk),
    .out(_U489_out)
);
assign _U490_in = in[4];
assign _U490_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U490 (
    .in(_U490_in),
    .clk(_U490_clk),
    .out(_U490_out)
);
assign out[4] = _U490_out;
assign out[3] = _U489_out;
assign out[2] = _U488_out;
assign out[1] = _U487_out;
assign out[0] = _U486_out;
endmodule

module array_delay_U478 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U479_in;
wire _U479_clk;
wire [15:0] _U479_out;
wire [15:0] _U480_in;
wire _U480_clk;
wire [15:0] _U480_out;
wire [15:0] _U481_in;
wire _U481_clk;
wire [15:0] _U481_out;
wire [15:0] _U482_in;
wire _U482_clk;
wire [15:0] _U482_out;
wire [15:0] _U483_in;
wire _U483_clk;
wire [15:0] _U483_out;
assign _U479_in = in[0];
assign _U479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(_U479_in),
    .clk(_U479_clk),
    .out(_U479_out)
);
assign _U480_in = in[1];
assign _U480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U480 (
    .in(_U480_in),
    .clk(_U480_clk),
    .out(_U480_out)
);
assign _U481_in = in[2];
assign _U481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U481_in),
    .clk(_U481_clk),
    .out(_U481_out)
);
assign _U482_in = in[3];
assign _U482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U482_in),
    .clk(_U482_clk),
    .out(_U482_out)
);
assign _U483_in = in[4];
assign _U483_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U483 (
    .in(_U483_in),
    .clk(_U483_clk),
    .out(_U483_out)
);
assign out[4] = _U483_out;
assign out[3] = _U482_out;
assign out[2] = _U481_out;
assign out[1] = _U480_out;
assign out[0] = _U479_out;
endmodule

module array_delay_U471 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U472_in;
wire _U472_clk;
wire [15:0] _U472_out;
wire [15:0] _U473_in;
wire _U473_clk;
wire [15:0] _U473_out;
wire [15:0] _U474_in;
wire _U474_clk;
wire [15:0] _U474_out;
wire [15:0] _U475_in;
wire _U475_clk;
wire [15:0] _U475_out;
wire [15:0] _U476_in;
wire _U476_clk;
wire [15:0] _U476_out;
assign _U472_in = in[0];
assign _U472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U472 (
    .in(_U472_in),
    .clk(_U472_clk),
    .out(_U472_out)
);
assign _U473_in = in[1];
assign _U473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U473 (
    .in(_U473_in),
    .clk(_U473_clk),
    .out(_U473_out)
);
assign _U474_in = in[2];
assign _U474_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U474 (
    .in(_U474_in),
    .clk(_U474_clk),
    .out(_U474_out)
);
assign _U475_in = in[3];
assign _U475_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U475 (
    .in(_U475_in),
    .clk(_U475_clk),
    .out(_U475_out)
);
assign _U476_in = in[4];
assign _U476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(_U476_in),
    .clk(_U476_clk),
    .out(_U476_out)
);
assign out[4] = _U476_out;
assign out[3] = _U475_out;
assign out[2] = _U474_out;
assign out[1] = _U473_out;
assign out[0] = _U472_out;
endmodule

module array_delay_U464 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire _U466_clk;
wire [15:0] _U466_out;
wire [15:0] _U467_in;
wire _U467_clk;
wire [15:0] _U467_out;
wire [15:0] _U468_in;
wire _U468_clk;
wire [15:0] _U468_out;
wire [15:0] _U469_in;
wire _U469_clk;
wire [15:0] _U469_out;
assign _U465_in = in[0];
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = in[1];
assign _U466_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U466 (
    .in(_U466_in),
    .clk(_U466_clk),
    .out(_U466_out)
);
assign _U467_in = in[2];
assign _U467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U467 (
    .in(_U467_in),
    .clk(_U467_clk),
    .out(_U467_out)
);
assign _U468_in = in[3];
assign _U468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U468_in),
    .clk(_U468_clk),
    .out(_U468_out)
);
assign _U469_in = in[4];
assign _U469_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U469 (
    .in(_U469_in),
    .clk(_U469_clk),
    .out(_U469_out)
);
assign out[4] = _U469_out;
assign out[3] = _U468_out;
assign out[2] = _U467_out;
assign out[1] = _U466_out;
assign out[0] = _U465_out;
endmodule

module array_delay_U457 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U458_in;
wire _U458_clk;
wire [15:0] _U458_out;
wire [15:0] _U459_in;
wire _U459_clk;
wire [15:0] _U459_out;
wire [15:0] _U460_in;
wire _U460_clk;
wire [15:0] _U460_out;
wire [15:0] _U461_in;
wire _U461_clk;
wire [15:0] _U461_out;
wire [15:0] _U462_in;
wire _U462_clk;
wire [15:0] _U462_out;
assign _U458_in = in[0];
assign _U458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U458 (
    .in(_U458_in),
    .clk(_U458_clk),
    .out(_U458_out)
);
assign _U459_in = in[1];
assign _U459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U459 (
    .in(_U459_in),
    .clk(_U459_clk),
    .out(_U459_out)
);
assign _U460_in = in[2];
assign _U460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U460 (
    .in(_U460_in),
    .clk(_U460_clk),
    .out(_U460_out)
);
assign _U461_in = in[3];
assign _U461_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U461 (
    .in(_U461_in),
    .clk(_U461_clk),
    .out(_U461_out)
);
assign _U462_in = in[4];
assign _U462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U462_in),
    .clk(_U462_clk),
    .out(_U462_out)
);
assign out[4] = _U462_out;
assign out[3] = _U461_out;
assign out[2] = _U460_out;
assign out[1] = _U459_out;
assign out[0] = _U458_out;
endmodule

module array_delay_U450 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U451_in;
wire _U451_clk;
wire [15:0] _U451_out;
wire [15:0] _U452_in;
wire _U452_clk;
wire [15:0] _U452_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
wire [15:0] _U454_in;
wire _U454_clk;
wire [15:0] _U454_out;
wire [15:0] _U455_in;
wire _U455_clk;
wire [15:0] _U455_out;
assign _U451_in = in[0];
assign _U451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(_U451_in),
    .clk(_U451_clk),
    .out(_U451_out)
);
assign _U452_in = in[1];
assign _U452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U452_in),
    .clk(_U452_clk),
    .out(_U452_out)
);
assign _U453_in = in[2];
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign _U454_in = in[3];
assign _U454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U454 (
    .in(_U454_in),
    .clk(_U454_clk),
    .out(_U454_out)
);
assign _U455_in = in[4];
assign _U455_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U455 (
    .in(_U455_in),
    .clk(_U455_clk),
    .out(_U455_out)
);
assign out[4] = _U455_out;
assign out[3] = _U454_out;
assign out[2] = _U453_out;
assign out[1] = _U452_out;
assign out[0] = _U451_out;
endmodule

module array_delay_U45 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U46_in;
wire _U46_clk;
wire [15:0] _U46_out;
wire [15:0] _U47_in;
wire _U47_clk;
wire [15:0] _U47_out;
wire [15:0] _U48_in;
wire _U48_clk;
wire [15:0] _U48_out;
wire [15:0] _U49_in;
wire _U49_clk;
wire [15:0] _U49_out;
assign _U46_in = in[0];
assign _U46_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(_U46_in),
    .clk(_U46_clk),
    .out(_U46_out)
);
assign _U47_in = in[1];
assign _U47_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U47 (
    .in(_U47_in),
    .clk(_U47_clk),
    .out(_U47_out)
);
assign _U48_in = in[2];
assign _U48_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U48 (
    .in(_U48_in),
    .clk(_U48_clk),
    .out(_U48_out)
);
assign _U49_in = in[3];
assign _U49_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U49_in),
    .clk(_U49_clk),
    .out(_U49_out)
);
assign out[3] = _U49_out;
assign out[2] = _U48_out;
assign out[1] = _U47_out;
assign out[0] = _U46_out;
endmodule

module array_delay_U443 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
wire [15:0] _U447_in;
wire _U447_clk;
wire [15:0] _U447_out;
wire [15:0] _U448_in;
wire _U448_clk;
wire [15:0] _U448_out;
assign _U444_in = in[0];
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = in[1];
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = in[2];
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign _U447_in = in[3];
assign _U447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U447 (
    .in(_U447_in),
    .clk(_U447_clk),
    .out(_U447_out)
);
assign _U448_in = in[4];
assign _U448_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U448 (
    .in(_U448_in),
    .clk(_U448_clk),
    .out(_U448_out)
);
assign out[4] = _U448_out;
assign out[3] = _U447_out;
assign out[2] = _U446_out;
assign out[1] = _U445_out;
assign out[0] = _U444_out;
endmodule

module array_delay_U436 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U437_in;
wire _U437_clk;
wire [15:0] _U437_out;
wire [15:0] _U438_in;
wire _U438_clk;
wire [15:0] _U438_out;
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
assign _U437_in = in[0];
assign _U437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U437 (
    .in(_U437_in),
    .clk(_U437_clk),
    .out(_U437_out)
);
assign _U438_in = in[1];
assign _U438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(_U438_in),
    .clk(_U438_clk),
    .out(_U438_out)
);
assign _U439_in = in[2];
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign _U440_in = in[3];
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = in[4];
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign out[4] = _U441_out;
assign out[3] = _U440_out;
assign out[2] = _U439_out;
assign out[1] = _U438_out;
assign out[0] = _U437_out;
endmodule

module array_delay_U429 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U430_in;
wire _U430_clk;
wire [15:0] _U430_out;
wire [15:0] _U431_in;
wire _U431_clk;
wire [15:0] _U431_out;
wire [15:0] _U432_in;
wire _U432_clk;
wire [15:0] _U432_out;
wire [15:0] _U433_in;
wire _U433_clk;
wire [15:0] _U433_out;
wire [15:0] _U434_in;
wire _U434_clk;
wire [15:0] _U434_out;
assign _U430_in = in[0];
assign _U430_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U430 (
    .in(_U430_in),
    .clk(_U430_clk),
    .out(_U430_out)
);
assign _U431_in = in[1];
assign _U431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U431_in),
    .clk(_U431_clk),
    .out(_U431_out)
);
assign _U432_in = in[2];
assign _U432_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U432 (
    .in(_U432_in),
    .clk(_U432_clk),
    .out(_U432_out)
);
assign _U433_in = in[3];
assign _U433_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U433 (
    .in(_U433_in),
    .clk(_U433_clk),
    .out(_U433_out)
);
assign _U434_in = in[4];
assign _U434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U434_in),
    .clk(_U434_clk),
    .out(_U434_out)
);
assign out[4] = _U434_out;
assign out[3] = _U433_out;
assign out[2] = _U432_out;
assign out[1] = _U431_out;
assign out[0] = _U430_out;
endmodule

module array_delay_U403 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U404_in;
wire _U404_clk;
wire [15:0] _U404_out;
wire [15:0] _U405_in;
wire _U405_clk;
wire [15:0] _U405_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire _U407_clk;
wire [15:0] _U407_out;
wire [15:0] _U408_in;
wire _U408_clk;
wire [15:0] _U408_out;
assign _U404_in = in[0];
assign _U404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U404 (
    .in(_U404_in),
    .clk(_U404_clk),
    .out(_U404_out)
);
assign _U405_in = in[1];
assign _U405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(_U405_in),
    .clk(_U405_clk),
    .out(_U405_out)
);
assign _U406_in = in[2];
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = in[3];
assign _U407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U407 (
    .in(_U407_in),
    .clk(_U407_clk),
    .out(_U407_out)
);
assign _U408_in = in[4];
assign _U408_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U408 (
    .in(_U408_in),
    .clk(_U408_clk),
    .out(_U408_out)
);
assign out[4] = _U408_out;
assign out[3] = _U407_out;
assign out[2] = _U406_out;
assign out[1] = _U405_out;
assign out[0] = _U404_out;
endmodule

module array_delay_U396 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U397_in;
wire _U397_clk;
wire [15:0] _U397_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
wire [15:0] _U400_in;
wire _U400_clk;
wire [15:0] _U400_out;
wire [15:0] _U401_in;
wire _U401_clk;
wire [15:0] _U401_out;
assign _U397_in = in[0];
assign _U397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U397_in),
    .clk(_U397_clk),
    .out(_U397_out)
);
assign _U398_in = in[1];
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = in[2];
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign _U400_in = in[3];
assign _U400_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U400 (
    .in(_U400_in),
    .clk(_U400_clk),
    .out(_U400_out)
);
assign _U401_in = in[4];
assign _U401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U401_in),
    .clk(_U401_clk),
    .out(_U401_out)
);
assign out[4] = _U401_out;
assign out[3] = _U400_out;
assign out[2] = _U399_out;
assign out[1] = _U398_out;
assign out[0] = _U397_out;
endmodule

module array_delay_U375 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U376_in;
wire _U376_clk;
wire [15:0] _U376_out;
wire [15:0] _U377_in;
wire _U377_clk;
wire [15:0] _U377_out;
wire [15:0] _U378_in;
wire _U378_clk;
wire [15:0] _U378_out;
wire [15:0] _U379_in;
wire _U379_clk;
wire [15:0] _U379_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
assign _U376_in = in[0];
assign _U376_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U376 (
    .in(_U376_in),
    .clk(_U376_clk),
    .out(_U376_out)
);
assign _U377_in = in[1];
assign _U377_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U377 (
    .in(_U377_in),
    .clk(_U377_clk),
    .out(_U377_out)
);
assign _U378_in = in[2];
assign _U378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U378_in),
    .clk(_U378_clk),
    .out(_U378_out)
);
assign _U379_in = in[3];
assign _U379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U379_in),
    .clk(_U379_clk),
    .out(_U379_out)
);
assign _U380_in = in[4];
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign out[4] = _U380_out;
assign out[3] = _U379_out;
assign out[2] = _U378_out;
assign out[1] = _U377_out;
assign out[0] = _U376_out;
endmodule

module array_delay_U368 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U369_in;
wire _U369_clk;
wire [15:0] _U369_out;
wire [15:0] _U370_in;
wire _U370_clk;
wire [15:0] _U370_out;
wire [15:0] _U371_in;
wire _U371_clk;
wire [15:0] _U371_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire _U373_clk;
wire [15:0] _U373_out;
assign _U369_in = in[0];
assign _U369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U369 (
    .in(_U369_in),
    .clk(_U369_clk),
    .out(_U369_out)
);
assign _U370_in = in[1];
assign _U370_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U370 (
    .in(_U370_in),
    .clk(_U370_clk),
    .out(_U370_out)
);
assign _U371_in = in[2];
assign _U371_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(_U371_in),
    .clk(_U371_clk),
    .out(_U371_out)
);
assign _U372_in = in[3];
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = in[4];
assign _U373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U373 (
    .in(_U373_in),
    .clk(_U373_clk),
    .out(_U373_out)
);
assign out[4] = _U373_out;
assign out[3] = _U372_out;
assign out[2] = _U371_out;
assign out[1] = _U370_out;
assign out[0] = _U369_out;
endmodule

module array_delay_U361 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U362_in;
wire _U362_clk;
wire [15:0] _U362_out;
wire [15:0] _U363_in;
wire _U363_clk;
wire [15:0] _U363_out;
wire [15:0] _U364_in;
wire _U364_clk;
wire [15:0] _U364_out;
wire [15:0] _U365_in;
wire _U365_clk;
wire [15:0] _U365_out;
wire [15:0] _U366_in;
wire _U366_clk;
wire [15:0] _U366_out;
assign _U362_in = in[0];
assign _U362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U362 (
    .in(_U362_in),
    .clk(_U362_clk),
    .out(_U362_out)
);
assign _U363_in = in[1];
assign _U363_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U363 (
    .in(_U363_in),
    .clk(_U363_clk),
    .out(_U363_out)
);
assign _U364_in = in[2];
assign _U364_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U364 (
    .in(_U364_in),
    .clk(_U364_clk),
    .out(_U364_out)
);
assign _U365_in = in[3];
assign _U365_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U365 (
    .in(_U365_in),
    .clk(_U365_clk),
    .out(_U365_out)
);
assign _U366_in = in[4];
assign _U366_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U366 (
    .in(_U366_in),
    .clk(_U366_clk),
    .out(_U366_out)
);
assign out[4] = _U366_out;
assign out[3] = _U365_out;
assign out[2] = _U364_out;
assign out[1] = _U363_out;
assign out[0] = _U362_out;
endmodule

module array_delay_U354 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire _U356_clk;
wire [15:0] _U356_out;
wire [15:0] _U357_in;
wire _U357_clk;
wire [15:0] _U357_out;
wire [15:0] _U358_in;
wire _U358_clk;
wire [15:0] _U358_out;
wire [15:0] _U359_in;
wire _U359_clk;
wire [15:0] _U359_out;
assign _U355_in = in[0];
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = in[1];
assign _U356_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U356 (
    .in(_U356_in),
    .clk(_U356_clk),
    .out(_U356_out)
);
assign _U357_in = in[2];
assign _U357_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U357 (
    .in(_U357_in),
    .clk(_U357_clk),
    .out(_U357_out)
);
assign _U358_in = in[3];
assign _U358_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U358 (
    .in(_U358_in),
    .clk(_U358_clk),
    .out(_U358_out)
);
assign _U359_in = in[4];
assign _U359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U359 (
    .in(_U359_in),
    .clk(_U359_clk),
    .out(_U359_out)
);
assign out[4] = _U359_out;
assign out[3] = _U358_out;
assign out[2] = _U357_out;
assign out[1] = _U356_out;
assign out[0] = _U355_out;
endmodule

module array_delay_U35 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U36_in;
wire _U36_clk;
wire [15:0] _U36_out;
wire [15:0] _U37_in;
wire _U37_clk;
wire [15:0] _U37_out;
wire [15:0] _U38_in;
wire _U38_clk;
wire [15:0] _U38_out;
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
assign _U36_in = in[0];
assign _U36_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(_U36_in),
    .clk(_U36_clk),
    .out(_U36_out)
);
assign _U37_in = in[1];
assign _U37_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U37 (
    .in(_U37_in),
    .clk(_U37_clk),
    .out(_U37_out)
);
assign _U38_in = in[2];
assign _U38_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U38 (
    .in(_U38_in),
    .clk(_U38_clk),
    .out(_U38_out)
);
assign _U39_in = in[3];
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign out[3] = _U39_out;
assign out[2] = _U38_out;
assign out[1] = _U37_out;
assign out[0] = _U36_out;
endmodule

module array_delay_U347 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U348_in;
wire _U348_clk;
wire [15:0] _U348_out;
wire [15:0] _U349_in;
wire _U349_clk;
wire [15:0] _U349_out;
wire [15:0] _U350_in;
wire _U350_clk;
wire [15:0] _U350_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire _U352_clk;
wire [15:0] _U352_out;
assign _U348_in = in[0];
assign _U348_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U348 (
    .in(_U348_in),
    .clk(_U348_clk),
    .out(_U348_out)
);
assign _U349_in = in[1];
assign _U349_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U349 (
    .in(_U349_in),
    .clk(_U349_clk),
    .out(_U349_out)
);
assign _U350_in = in[2];
assign _U350_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U350_in),
    .clk(_U350_clk),
    .out(_U350_out)
);
assign _U351_in = in[3];
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = in[4];
assign _U352_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U352 (
    .in(_U352_in),
    .clk(_U352_clk),
    .out(_U352_out)
);
assign out[4] = _U352_out;
assign out[3] = _U351_out;
assign out[2] = _U350_out;
assign out[1] = _U349_out;
assign out[0] = _U348_out;
endmodule

module array_delay_U340 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire _U342_clk;
wire [15:0] _U342_out;
wire [15:0] _U343_in;
wire _U343_clk;
wire [15:0] _U343_out;
wire [15:0] _U344_in;
wire _U344_clk;
wire [15:0] _U344_out;
wire [15:0] _U345_in;
wire _U345_clk;
wire [15:0] _U345_out;
assign _U341_in = in[0];
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = in[1];
assign _U342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U342_in),
    .clk(_U342_clk),
    .out(_U342_out)
);
assign _U343_in = in[2];
assign _U343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U343 (
    .in(_U343_in),
    .clk(_U343_clk),
    .out(_U343_out)
);
assign _U344_in = in[3];
assign _U344_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U344 (
    .in(_U344_in),
    .clk(_U344_clk),
    .out(_U344_out)
);
assign _U345_in = in[4];
assign _U345_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(_U345_in),
    .clk(_U345_clk),
    .out(_U345_out)
);
assign out[4] = _U345_out;
assign out[3] = _U344_out;
assign out[2] = _U343_out;
assign out[1] = _U342_out;
assign out[0] = _U341_out;
endmodule

module array_delay_U333 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U334_in;
wire _U334_clk;
wire [15:0] _U334_out;
wire [15:0] _U335_in;
wire _U335_clk;
wire [15:0] _U335_out;
wire [15:0] _U336_in;
wire _U336_clk;
wire [15:0] _U336_out;
wire [15:0] _U337_in;
wire _U337_clk;
wire [15:0] _U337_out;
wire [15:0] _U338_in;
wire _U338_clk;
wire [15:0] _U338_out;
assign _U334_in = in[0];
assign _U334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U334 (
    .in(_U334_in),
    .clk(_U334_clk),
    .out(_U334_out)
);
assign _U335_in = in[1];
assign _U335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U335 (
    .in(_U335_in),
    .clk(_U335_clk),
    .out(_U335_out)
);
assign _U336_in = in[2];
assign _U336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(_U336_in),
    .clk(_U336_clk),
    .out(_U336_out)
);
assign _U337_in = in[3];
assign _U337_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U337 (
    .in(_U337_in),
    .clk(_U337_clk),
    .out(_U337_out)
);
assign _U338_in = in[4];
assign _U338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U338_in),
    .clk(_U338_clk),
    .out(_U338_out)
);
assign out[4] = _U338_out;
assign out[3] = _U337_out;
assign out[2] = _U336_out;
assign out[1] = _U335_out;
assign out[0] = _U334_out;
endmodule

module array_delay_U326 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U327_in;
wire _U327_clk;
wire [15:0] _U327_out;
wire [15:0] _U328_in;
wire _U328_clk;
wire [15:0] _U328_out;
wire [15:0] _U329_in;
wire _U329_clk;
wire [15:0] _U329_out;
wire [15:0] _U330_in;
wire _U330_clk;
wire [15:0] _U330_out;
wire [15:0] _U331_in;
wire _U331_clk;
wire [15:0] _U331_out;
assign _U327_in = in[0];
assign _U327_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U327 (
    .in(_U327_in),
    .clk(_U327_clk),
    .out(_U327_out)
);
assign _U328_in = in[1];
assign _U328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U328_in),
    .clk(_U328_clk),
    .out(_U328_out)
);
assign _U329_in = in[2];
assign _U329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U329 (
    .in(_U329_in),
    .clk(_U329_clk),
    .out(_U329_out)
);
assign _U330_in = in[3];
assign _U330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U330_in),
    .clk(_U330_clk),
    .out(_U330_out)
);
assign _U331_in = in[4];
assign _U331_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U331 (
    .in(_U331_in),
    .clk(_U331_clk),
    .out(_U331_out)
);
assign out[4] = _U331_out;
assign out[3] = _U330_out;
assign out[2] = _U329_out;
assign out[1] = _U328_out;
assign out[0] = _U327_out;
endmodule

module array_delay_U319 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U320_in;
wire _U320_clk;
wire [15:0] _U320_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire _U322_clk;
wire [15:0] _U322_out;
wire [15:0] _U323_in;
wire _U323_clk;
wire [15:0] _U323_out;
wire [15:0] _U324_in;
wire _U324_clk;
wire [15:0] _U324_out;
assign _U320_in = in[0];
assign _U320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U320_in),
    .clk(_U320_clk),
    .out(_U320_out)
);
assign _U321_in = in[1];
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = in[2];
assign _U322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U322 (
    .in(_U322_in),
    .clk(_U322_clk),
    .out(_U322_out)
);
assign _U323_in = in[3];
assign _U323_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U323 (
    .in(_U323_in),
    .clk(_U323_clk),
    .out(_U323_out)
);
assign _U324_in = in[4];
assign _U324_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U324 (
    .in(_U324_in),
    .clk(_U324_clk),
    .out(_U324_out)
);
assign out[4] = _U324_out;
assign out[3] = _U323_out;
assign out[2] = _U322_out;
assign out[1] = _U321_out;
assign out[0] = _U320_out;
endmodule

module array_delay_U312 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U313_in;
wire _U313_clk;
wire [15:0] _U313_out;
wire [15:0] _U314_in;
wire _U314_clk;
wire [15:0] _U314_out;
wire [15:0] _U315_in;
wire _U315_clk;
wire [15:0] _U315_out;
wire [15:0] _U316_in;
wire _U316_clk;
wire [15:0] _U316_out;
wire [15:0] _U317_in;
wire _U317_clk;
wire [15:0] _U317_out;
assign _U313_in = in[0];
assign _U313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U313 (
    .in(_U313_in),
    .clk(_U313_clk),
    .out(_U313_out)
);
assign _U314_in = in[1];
assign _U314_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U314 (
    .in(_U314_in),
    .clk(_U314_clk),
    .out(_U314_out)
);
assign _U315_in = in[2];
assign _U315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U315_in),
    .clk(_U315_clk),
    .out(_U315_out)
);
assign _U316_in = in[3];
assign _U316_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U316 (
    .in(_U316_in),
    .clk(_U316_clk),
    .out(_U316_out)
);
assign _U317_in = in[4];
assign _U317_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U317 (
    .in(_U317_in),
    .clk(_U317_clk),
    .out(_U317_out)
);
assign out[4] = _U317_out;
assign out[3] = _U316_out;
assign out[2] = _U315_out;
assign out[1] = _U314_out;
assign out[0] = _U313_out;
endmodule

module array_delay_U305 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U306_in;
wire _U306_clk;
wire [15:0] _U306_out;
wire [15:0] _U307_in;
wire _U307_clk;
wire [15:0] _U307_out;
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire _U310_clk;
wire [15:0] _U310_out;
assign _U306_in = in[0];
assign _U306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U306_in),
    .clk(_U306_clk),
    .out(_U306_out)
);
assign _U307_in = in[1];
assign _U307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U307 (
    .in(_U307_in),
    .clk(_U307_clk),
    .out(_U307_out)
);
assign _U308_in = in[2];
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = in[3];
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = in[4];
assign _U310_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U310 (
    .in(_U310_in),
    .clk(_U310_clk),
    .out(_U310_out)
);
assign out[4] = _U310_out;
assign out[3] = _U309_out;
assign out[2] = _U308_out;
assign out[1] = _U307_out;
assign out[0] = _U306_out;
endmodule

module array_delay_U298 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U299_in;
wire _U299_clk;
wire [15:0] _U299_out;
wire [15:0] _U300_in;
wire _U300_clk;
wire [15:0] _U300_out;
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire _U303_clk;
wire [15:0] _U303_out;
assign _U299_in = in[0];
assign _U299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U299_in),
    .clk(_U299_clk),
    .out(_U299_out)
);
assign _U300_in = in[1];
assign _U300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U300 (
    .in(_U300_in),
    .clk(_U300_clk),
    .out(_U300_out)
);
assign _U301_in = in[2];
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = in[3];
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = in[4];
assign _U303_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U303 (
    .in(_U303_in),
    .clk(_U303_clk),
    .out(_U303_out)
);
assign out[4] = _U303_out;
assign out[3] = _U302_out;
assign out[2] = _U301_out;
assign out[1] = _U300_out;
assign out[0] = _U299_out;
endmodule

module array_delay_U291 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U292_in;
wire _U292_clk;
wire [15:0] _U292_out;
wire [15:0] _U293_in;
wire _U293_clk;
wire [15:0] _U293_out;
wire [15:0] _U294_in;
wire _U294_clk;
wire [15:0] _U294_out;
wire [15:0] _U295_in;
wire _U295_clk;
wire [15:0] _U295_out;
wire [15:0] _U296_in;
wire _U296_clk;
wire [15:0] _U296_out;
assign _U292_in = in[0];
assign _U292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U292 (
    .in(_U292_in),
    .clk(_U292_clk),
    .out(_U292_out)
);
assign _U293_in = in[1];
assign _U293_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U293 (
    .in(_U293_in),
    .clk(_U293_clk),
    .out(_U293_out)
);
assign _U294_in = in[2];
assign _U294_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U294 (
    .in(_U294_in),
    .clk(_U294_clk),
    .out(_U294_out)
);
assign _U295_in = in[3];
assign _U295_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U295 (
    .in(_U295_in),
    .clk(_U295_clk),
    .out(_U295_out)
);
assign _U296_in = in[4];
assign _U296_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U296 (
    .in(_U296_in),
    .clk(_U296_clk),
    .out(_U296_out)
);
assign out[4] = _U296_out;
assign out[3] = _U295_out;
assign out[2] = _U294_out;
assign out[1] = _U293_out;
assign out[0] = _U292_out;
endmodule

module array_delay_U29 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U30_in;
wire _U30_clk;
wire [15:0] _U30_out;
wire [15:0] _U31_in;
wire _U31_clk;
wire [15:0] _U31_out;
wire [15:0] _U32_in;
wire _U32_clk;
wire [15:0] _U32_out;
wire [15:0] _U33_in;
wire _U33_clk;
wire [15:0] _U33_out;
assign _U30_in = in[0];
assign _U30_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U30 (
    .in(_U30_in),
    .clk(_U30_clk),
    .out(_U30_out)
);
assign _U31_in = in[1];
assign _U31_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U31 (
    .in(_U31_in),
    .clk(_U31_clk),
    .out(_U31_out)
);
assign _U32_in = in[2];
assign _U32_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U32 (
    .in(_U32_in),
    .clk(_U32_clk),
    .out(_U32_out)
);
assign _U33_in = in[3];
assign _U33_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U33 (
    .in(_U33_in),
    .clk(_U33_clk),
    .out(_U33_out)
);
assign out[3] = _U33_out;
assign out[2] = _U32_out;
assign out[1] = _U31_out;
assign out[0] = _U30_out;
endmodule

module array_delay_U284 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U285_in;
wire _U285_clk;
wire [15:0] _U285_out;
wire [15:0] _U286_in;
wire _U286_clk;
wire [15:0] _U286_out;
wire [15:0] _U287_in;
wire _U287_clk;
wire [15:0] _U287_out;
wire [15:0] _U288_in;
wire _U288_clk;
wire [15:0] _U288_out;
wire [15:0] _U289_in;
wire _U289_clk;
wire [15:0] _U289_out;
assign _U285_in = in[0];
assign _U285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(_U285_in),
    .clk(_U285_clk),
    .out(_U285_out)
);
assign _U286_in = in[1];
assign _U286_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U286 (
    .in(_U286_in),
    .clk(_U286_clk),
    .out(_U286_out)
);
assign _U287_in = in[2];
assign _U287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U287 (
    .in(_U287_in),
    .clk(_U287_clk),
    .out(_U287_out)
);
assign _U288_in = in[3];
assign _U288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U288_in),
    .clk(_U288_clk),
    .out(_U288_out)
);
assign _U289_in = in[4];
assign _U289_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U289_in),
    .clk(_U289_clk),
    .out(_U289_out)
);
assign out[4] = _U289_out;
assign out[3] = _U288_out;
assign out[2] = _U287_out;
assign out[1] = _U286_out;
assign out[0] = _U285_out;
endmodule

module array_delay_U277 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire _U279_clk;
wire [15:0] _U279_out;
wire [15:0] _U280_in;
wire _U280_clk;
wire [15:0] _U280_out;
wire [15:0] _U281_in;
wire _U281_clk;
wire [15:0] _U281_out;
wire [15:0] _U282_in;
wire _U282_clk;
wire [15:0] _U282_out;
assign _U278_in = in[0];
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = in[1];
assign _U279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U279_in),
    .clk(_U279_clk),
    .out(_U279_out)
);
assign _U280_in = in[2];
assign _U280_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U280 (
    .in(_U280_in),
    .clk(_U280_clk),
    .out(_U280_out)
);
assign _U281_in = in[3];
assign _U281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U281_in),
    .clk(_U281_clk),
    .out(_U281_out)
);
assign _U282_in = in[4];
assign _U282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U282 (
    .in(_U282_in),
    .clk(_U282_clk),
    .out(_U282_out)
);
assign out[4] = _U282_out;
assign out[3] = _U281_out;
assign out[2] = _U280_out;
assign out[1] = _U279_out;
assign out[0] = _U278_out;
endmodule

module array_delay_U270 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U271_in;
wire _U271_clk;
wire [15:0] _U271_out;
wire [15:0] _U272_in;
wire _U272_clk;
wire [15:0] _U272_out;
wire [15:0] _U273_in;
wire _U273_clk;
wire [15:0] _U273_out;
wire [15:0] _U274_in;
wire _U274_clk;
wire [15:0] _U274_out;
wire [15:0] _U275_in;
wire _U275_clk;
wire [15:0] _U275_out;
assign _U271_in = in[0];
assign _U271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U271_in),
    .clk(_U271_clk),
    .out(_U271_out)
);
assign _U272_in = in[1];
assign _U272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U272_in),
    .clk(_U272_clk),
    .out(_U272_out)
);
assign _U273_in = in[2];
assign _U273_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U273 (
    .in(_U273_in),
    .clk(_U273_clk),
    .out(_U273_out)
);
assign _U274_in = in[3];
assign _U274_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U274 (
    .in(_U274_in),
    .clk(_U274_clk),
    .out(_U274_out)
);
assign _U275_in = in[4];
assign _U275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U275 (
    .in(_U275_in),
    .clk(_U275_clk),
    .out(_U275_out)
);
assign out[4] = _U275_out;
assign out[3] = _U274_out;
assign out[2] = _U273_out;
assign out[1] = _U272_out;
assign out[0] = _U271_out;
endmodule

module array_delay_U263 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U264_in;
wire _U264_clk;
wire [15:0] _U264_out;
wire [15:0] _U265_in;
wire _U265_clk;
wire [15:0] _U265_out;
wire [15:0] _U266_in;
wire _U266_clk;
wire [15:0] _U266_out;
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire _U268_clk;
wire [15:0] _U268_out;
assign _U264_in = in[0];
assign _U264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U264_in),
    .clk(_U264_clk),
    .out(_U264_out)
);
assign _U265_in = in[1];
assign _U265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U265 (
    .in(_U265_in),
    .clk(_U265_clk),
    .out(_U265_out)
);
assign _U266_in = in[2];
assign _U266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U266 (
    .in(_U266_in),
    .clk(_U266_clk),
    .out(_U266_out)
);
assign _U267_in = in[3];
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = in[4];
assign _U268_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U268 (
    .in(_U268_in),
    .clk(_U268_clk),
    .out(_U268_out)
);
assign out[4] = _U268_out;
assign out[3] = _U267_out;
assign out[2] = _U266_out;
assign out[1] = _U265_out;
assign out[0] = _U264_out;
endmodule

module array_delay_U237 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U238_in;
wire _U238_clk;
wire [15:0] _U238_out;
wire [15:0] _U239_in;
wire _U239_clk;
wire [15:0] _U239_out;
wire [15:0] _U240_in;
wire _U240_clk;
wire [15:0] _U240_out;
wire [15:0] _U241_in;
wire _U241_clk;
wire [15:0] _U241_out;
wire [15:0] _U242_in;
wire _U242_clk;
wire [15:0] _U242_out;
assign _U238_in = in[0];
assign _U238_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U238 (
    .in(_U238_in),
    .clk(_U238_clk),
    .out(_U238_out)
);
assign _U239_in = in[1];
assign _U239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U239 (
    .in(_U239_in),
    .clk(_U239_clk),
    .out(_U239_out)
);
assign _U240_in = in[2];
assign _U240_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U240 (
    .in(_U240_in),
    .clk(_U240_clk),
    .out(_U240_out)
);
assign _U241_in = in[3];
assign _U241_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U241 (
    .in(_U241_in),
    .clk(_U241_clk),
    .out(_U241_out)
);
assign _U242_in = in[4];
assign _U242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U242_in),
    .clk(_U242_clk),
    .out(_U242_out)
);
assign out[4] = _U242_out;
assign out[3] = _U241_out;
assign out[2] = _U240_out;
assign out[1] = _U239_out;
assign out[0] = _U238_out;
endmodule

module array_delay_U230 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U231_in;
wire _U231_clk;
wire [15:0] _U231_out;
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
wire [15:0] _U233_in;
wire _U233_clk;
wire [15:0] _U233_out;
wire [15:0] _U234_in;
wire _U234_clk;
wire [15:0] _U234_out;
wire [15:0] _U235_in;
wire _U235_clk;
wire [15:0] _U235_out;
assign _U231_in = in[0];
assign _U231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U231 (
    .in(_U231_in),
    .clk(_U231_clk),
    .out(_U231_out)
);
assign _U232_in = in[1];
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign _U233_in = in[2];
assign _U233_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U233 (
    .in(_U233_in),
    .clk(_U233_clk),
    .out(_U233_out)
);
assign _U234_in = in[3];
assign _U234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U234 (
    .in(_U234_in),
    .clk(_U234_clk),
    .out(_U234_out)
);
assign _U235_in = in[4];
assign _U235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U235 (
    .in(_U235_in),
    .clk(_U235_clk),
    .out(_U235_out)
);
assign out[4] = _U235_out;
assign out[3] = _U234_out;
assign out[2] = _U233_out;
assign out[1] = _U232_out;
assign out[0] = _U231_out;
endmodule

module array_delay_U216 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
wire [15:0] _U219_in;
wire _U219_clk;
wire [15:0] _U219_out;
wire [15:0] _U220_in;
wire _U220_clk;
wire [15:0] _U220_out;
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
assign _U217_in = in[0];
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = in[1];
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign _U219_in = in[2];
assign _U219_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U219_in),
    .clk(_U219_clk),
    .out(_U219_out)
);
assign _U220_in = in[3];
assign _U220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U220_in),
    .clk(_U220_clk),
    .out(_U220_out)
);
assign _U221_in = in[4];
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign out[4] = _U221_out;
assign out[3] = _U220_out;
assign out[2] = _U219_out;
assign out[1] = _U218_out;
assign out[0] = _U217_out;
endmodule

module array_delay_U209 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U210_in;
wire _U210_clk;
wire [15:0] _U210_out;
wire [15:0] _U211_in;
wire _U211_clk;
wire [15:0] _U211_out;
wire [15:0] _U212_in;
wire _U212_clk;
wire [15:0] _U212_out;
wire [15:0] _U213_in;
wire _U213_clk;
wire [15:0] _U213_out;
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
assign _U210_in = in[0];
assign _U210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U210 (
    .in(_U210_in),
    .clk(_U210_clk),
    .out(_U210_out)
);
assign _U211_in = in[1];
assign _U211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(_U211_in),
    .clk(_U211_clk),
    .out(_U211_out)
);
assign _U212_in = in[2];
assign _U212_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U212 (
    .in(_U212_in),
    .clk(_U212_clk),
    .out(_U212_out)
);
assign _U213_in = in[3];
assign _U213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(_U213_in),
    .clk(_U213_clk),
    .out(_U213_out)
);
assign _U214_in = in[4];
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign out[4] = _U214_out;
assign out[3] = _U213_out;
assign out[2] = _U212_out;
assign out[1] = _U211_out;
assign out[0] = _U210_out;
endmodule

module array_delay_U202 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U203_in;
wire _U203_clk;
wire [15:0] _U203_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U205_in;
wire _U205_clk;
wire [15:0] _U205_out;
wire [15:0] _U206_in;
wire _U206_clk;
wire [15:0] _U206_out;
wire [15:0] _U207_in;
wire _U207_clk;
wire [15:0] _U207_out;
assign _U203_in = in[0];
assign _U203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U203 (
    .in(_U203_in),
    .clk(_U203_clk),
    .out(_U203_out)
);
assign _U204_in = in[1];
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U205_in = in[2];
assign _U205_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U205 (
    .in(_U205_in),
    .clk(_U205_clk),
    .out(_U205_out)
);
assign _U206_in = in[3];
assign _U206_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U206 (
    .in(_U206_in),
    .clk(_U206_clk),
    .out(_U206_out)
);
assign _U207_in = in[4];
assign _U207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(_U207_in),
    .clk(_U207_clk),
    .out(_U207_out)
);
assign out[4] = _U207_out;
assign out[3] = _U206_out;
assign out[2] = _U205_out;
assign out[1] = _U204_out;
assign out[0] = _U203_out;
endmodule

module array_delay_U195 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U196_in;
wire _U196_clk;
wire [15:0] _U196_out;
wire [15:0] _U197_in;
wire _U197_clk;
wire [15:0] _U197_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire _U199_clk;
wire [15:0] _U199_out;
wire [15:0] _U200_in;
wire _U200_clk;
wire [15:0] _U200_out;
assign _U196_in = in[0];
assign _U196_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U196 (
    .in(_U196_in),
    .clk(_U196_clk),
    .out(_U196_out)
);
assign _U197_in = in[1];
assign _U197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U197 (
    .in(_U197_in),
    .clk(_U197_clk),
    .out(_U197_out)
);
assign _U198_in = in[2];
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = in[3];
assign _U199_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U199 (
    .in(_U199_in),
    .clk(_U199_clk),
    .out(_U199_out)
);
assign _U200_in = in[4];
assign _U200_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U200 (
    .in(_U200_in),
    .clk(_U200_clk),
    .out(_U200_out)
);
assign out[4] = _U200_out;
assign out[3] = _U199_out;
assign out[2] = _U198_out;
assign out[1] = _U197_out;
assign out[0] = _U196_out;
endmodule

module array_delay_U188 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U189_in;
wire _U189_clk;
wire [15:0] _U189_out;
wire [15:0] _U190_in;
wire _U190_clk;
wire [15:0] _U190_out;
wire [15:0] _U191_in;
wire _U191_clk;
wire [15:0] _U191_out;
wire [15:0] _U192_in;
wire _U192_clk;
wire [15:0] _U192_out;
wire [15:0] _U193_in;
wire _U193_clk;
wire [15:0] _U193_out;
assign _U189_in = in[0];
assign _U189_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U189 (
    .in(_U189_in),
    .clk(_U189_clk),
    .out(_U189_out)
);
assign _U190_in = in[1];
assign _U190_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U190 (
    .in(_U190_in),
    .clk(_U190_clk),
    .out(_U190_out)
);
assign _U191_in = in[2];
assign _U191_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U191_in),
    .clk(_U191_clk),
    .out(_U191_out)
);
assign _U192_in = in[3];
assign _U192_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U192_in),
    .clk(_U192_clk),
    .out(_U192_out)
);
assign _U193_in = in[4];
assign _U193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U193_in),
    .clk(_U193_clk),
    .out(_U193_out)
);
assign out[4] = _U193_out;
assign out[3] = _U192_out;
assign out[2] = _U191_out;
assign out[1] = _U190_out;
assign out[0] = _U189_out;
endmodule

module array_delay_U181 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U182_in;
wire _U182_clk;
wire [15:0] _U182_out;
wire [15:0] _U183_in;
wire _U183_clk;
wire [15:0] _U183_out;
wire [15:0] _U184_in;
wire _U184_clk;
wire [15:0] _U184_out;
wire [15:0] _U185_in;
wire _U185_clk;
wire [15:0] _U185_out;
wire [15:0] _U186_in;
wire _U186_clk;
wire [15:0] _U186_out;
assign _U182_in = in[0];
assign _U182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U182_in),
    .clk(_U182_clk),
    .out(_U182_out)
);
assign _U183_in = in[1];
assign _U183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U183_in),
    .clk(_U183_clk),
    .out(_U183_out)
);
assign _U184_in = in[2];
assign _U184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U184_in),
    .clk(_U184_clk),
    .out(_U184_out)
);
assign _U185_in = in[3];
assign _U185_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U185 (
    .in(_U185_in),
    .clk(_U185_clk),
    .out(_U185_out)
);
assign _U186_in = in[4];
assign _U186_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U186 (
    .in(_U186_in),
    .clk(_U186_clk),
    .out(_U186_out)
);
assign out[4] = _U186_out;
assign out[3] = _U185_out;
assign out[2] = _U184_out;
assign out[1] = _U183_out;
assign out[0] = _U182_out;
endmodule

module array_delay_U174 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
wire [15:0] _U176_in;
wire _U176_clk;
wire [15:0] _U176_out;
wire [15:0] _U177_in;
wire _U177_clk;
wire [15:0] _U177_out;
wire [15:0] _U178_in;
wire _U178_clk;
wire [15:0] _U178_out;
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
assign _U175_in = in[0];
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign _U176_in = in[1];
assign _U176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U176 (
    .in(_U176_in),
    .clk(_U176_clk),
    .out(_U176_out)
);
assign _U177_in = in[2];
assign _U177_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U177 (
    .in(_U177_in),
    .clk(_U177_clk),
    .out(_U177_out)
);
assign _U178_in = in[3];
assign _U178_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U178 (
    .in(_U178_in),
    .clk(_U178_clk),
    .out(_U178_out)
);
assign _U179_in = in[4];
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign out[4] = _U179_out;
assign out[3] = _U178_out;
assign out[2] = _U177_out;
assign out[1] = _U176_out;
assign out[0] = _U175_out;
endmodule

module array_delay_U167 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
wire [15:0] _U169_in;
wire _U169_clk;
wire [15:0] _U169_out;
wire [15:0] _U170_in;
wire _U170_clk;
wire [15:0] _U170_out;
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire _U172_clk;
wire [15:0] _U172_out;
assign _U168_in = in[0];
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign _U169_in = in[1];
assign _U169_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U169 (
    .in(_U169_in),
    .clk(_U169_clk),
    .out(_U169_out)
);
assign _U170_in = in[2];
assign _U170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U170 (
    .in(_U170_in),
    .clk(_U170_clk),
    .out(_U170_out)
);
assign _U171_in = in[3];
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = in[4];
assign _U172_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(_U172_in),
    .clk(_U172_clk),
    .out(_U172_out)
);
assign out[4] = _U172_out;
assign out[3] = _U171_out;
assign out[2] = _U170_out;
assign out[1] = _U169_out;
assign out[0] = _U168_out;
endmodule

module array_delay_U160 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U161_in;
wire _U161_clk;
wire [15:0] _U161_out;
wire [15:0] _U162_in;
wire _U162_clk;
wire [15:0] _U162_out;
wire [15:0] _U163_in;
wire _U163_clk;
wire [15:0] _U163_out;
wire [15:0] _U164_in;
wire _U164_clk;
wire [15:0] _U164_out;
wire [15:0] _U165_in;
wire _U165_clk;
wire [15:0] _U165_out;
assign _U161_in = in[0];
assign _U161_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U161 (
    .in(_U161_in),
    .clk(_U161_clk),
    .out(_U161_out)
);
assign _U162_in = in[1];
assign _U162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(_U162_in),
    .clk(_U162_clk),
    .out(_U162_out)
);
assign _U163_in = in[2];
assign _U163_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(_U163_in),
    .clk(_U163_clk),
    .out(_U163_out)
);
assign _U164_in = in[3];
assign _U164_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(_U164_in),
    .clk(_U164_clk),
    .out(_U164_out)
);
assign _U165_in = in[4];
assign _U165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(_U165_in),
    .clk(_U165_clk),
    .out(_U165_out)
);
assign out[4] = _U165_out;
assign out[3] = _U164_out;
assign out[2] = _U163_out;
assign out[1] = _U162_out;
assign out[0] = _U161_out;
endmodule

module array_delay_U153 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U154_in;
wire _U154_clk;
wire [15:0] _U154_out;
wire [15:0] _U155_in;
wire _U155_clk;
wire [15:0] _U155_out;
wire [15:0] _U156_in;
wire _U156_clk;
wire [15:0] _U156_out;
wire [15:0] _U157_in;
wire _U157_clk;
wire [15:0] _U157_out;
wire [15:0] _U158_in;
wire _U158_clk;
wire [15:0] _U158_out;
assign _U154_in = in[0];
assign _U154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(_U154_in),
    .clk(_U154_clk),
    .out(_U154_out)
);
assign _U155_in = in[1];
assign _U155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U155_in),
    .clk(_U155_clk),
    .out(_U155_out)
);
assign _U156_in = in[2];
assign _U156_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U156 (
    .in(_U156_in),
    .clk(_U156_clk),
    .out(_U156_out)
);
assign _U157_in = in[3];
assign _U157_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U157 (
    .in(_U157_in),
    .clk(_U157_clk),
    .out(_U157_out)
);
assign _U158_in = in[4];
assign _U158_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U158 (
    .in(_U158_in),
    .clk(_U158_clk),
    .out(_U158_out)
);
assign out[4] = _U158_out;
assign out[3] = _U157_out;
assign out[2] = _U156_out;
assign out[1] = _U155_out;
assign out[0] = _U154_out;
endmodule

module array_delay_U146 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire _U148_clk;
wire [15:0] _U148_out;
wire [15:0] _U149_in;
wire _U149_clk;
wire [15:0] _U149_out;
wire [15:0] _U150_in;
wire _U150_clk;
wire [15:0] _U150_out;
wire [15:0] _U151_in;
wire _U151_clk;
wire [15:0] _U151_out;
assign _U147_in = in[0];
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = in[1];
assign _U148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U148_in),
    .clk(_U148_clk),
    .out(_U148_out)
);
assign _U149_in = in[2];
assign _U149_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U149 (
    .in(_U149_in),
    .clk(_U149_clk),
    .out(_U149_out)
);
assign _U150_in = in[3];
assign _U150_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U150 (
    .in(_U150_in),
    .clk(_U150_clk),
    .out(_U150_out)
);
assign _U151_in = in[4];
assign _U151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(_U151_in),
    .clk(_U151_clk),
    .out(_U151_out)
);
assign out[4] = _U151_out;
assign out[3] = _U150_out;
assign out[2] = _U149_out;
assign out[1] = _U148_out;
assign out[0] = _U147_out;
endmodule

module array_delay_U139 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire _U141_clk;
wire [15:0] _U141_out;
wire [15:0] _U142_in;
wire _U142_clk;
wire [15:0] _U142_out;
wire [15:0] _U143_in;
wire _U143_clk;
wire [15:0] _U143_out;
wire [15:0] _U144_in;
wire _U144_clk;
wire [15:0] _U144_out;
assign _U140_in = in[0];
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = in[1];
assign _U141_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U141 (
    .in(_U141_in),
    .clk(_U141_clk),
    .out(_U141_out)
);
assign _U142_in = in[2];
assign _U142_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U142 (
    .in(_U142_in),
    .clk(_U142_clk),
    .out(_U142_out)
);
assign _U143_in = in[3];
assign _U143_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U143 (
    .in(_U143_in),
    .clk(_U143_clk),
    .out(_U143_out)
);
assign _U144_in = in[4];
assign _U144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U144 (
    .in(_U144_in),
    .clk(_U144_clk),
    .out(_U144_out)
);
assign out[4] = _U144_out;
assign out[3] = _U143_out;
assign out[2] = _U142_out;
assign out[1] = _U141_out;
assign out[0] = _U140_out;
endmodule

module array_delay_U132 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U133_in;
wire _U133_clk;
wire [15:0] _U133_out;
wire [15:0] _U134_in;
wire _U134_clk;
wire [15:0] _U134_out;
wire [15:0] _U135_in;
wire _U135_clk;
wire [15:0] _U135_out;
wire [15:0] _U136_in;
wire _U136_clk;
wire [15:0] _U136_out;
wire [15:0] _U137_in;
wire _U137_clk;
wire [15:0] _U137_out;
assign _U133_in = in[0];
assign _U133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U133_in),
    .clk(_U133_clk),
    .out(_U133_out)
);
assign _U134_in = in[1];
assign _U134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U134_in),
    .clk(_U134_clk),
    .out(_U134_out)
);
assign _U135_in = in[2];
assign _U135_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U135 (
    .in(_U135_in),
    .clk(_U135_clk),
    .out(_U135_out)
);
assign _U136_in = in[3];
assign _U136_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U136 (
    .in(_U136_in),
    .clk(_U136_clk),
    .out(_U136_out)
);
assign _U137_in = in[4];
assign _U137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U137 (
    .in(_U137_in),
    .clk(_U137_clk),
    .out(_U137_out)
);
assign out[4] = _U137_out;
assign out[3] = _U136_out;
assign out[2] = _U135_out;
assign out[1] = _U134_out;
assign out[0] = _U133_out;
endmodule

module array_delay_U125 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U126_in;
wire _U126_clk;
wire [15:0] _U126_out;
wire [15:0] _U127_in;
wire _U127_clk;
wire [15:0] _U127_out;
wire [15:0] _U128_in;
wire _U128_clk;
wire [15:0] _U128_out;
wire [15:0] _U129_in;
wire _U129_clk;
wire [15:0] _U129_out;
wire [15:0] _U130_in;
wire _U130_clk;
wire [15:0] _U130_out;
assign _U126_in = in[0];
assign _U126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(_U126_in),
    .clk(_U126_clk),
    .out(_U126_out)
);
assign _U127_in = in[1];
assign _U127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U127_in),
    .clk(_U127_clk),
    .out(_U127_out)
);
assign _U128_in = in[2];
assign _U128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U128_in),
    .clk(_U128_clk),
    .out(_U128_out)
);
assign _U129_in = in[3];
assign _U129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U129_in),
    .clk(_U129_clk),
    .out(_U129_out)
);
assign _U130_in = in[4];
assign _U130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U130_in),
    .clk(_U130_clk),
    .out(_U130_out)
);
assign out[4] = _U130_out;
assign out[3] = _U129_out;
assign out[2] = _U128_out;
assign out[1] = _U127_out;
assign out[0] = _U126_out;
endmodule

module array_delay_U118 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U119_in;
wire _U119_clk;
wire [15:0] _U119_out;
wire [15:0] _U120_in;
wire _U120_clk;
wire [15:0] _U120_out;
wire [15:0] _U121_in;
wire _U121_clk;
wire [15:0] _U121_out;
wire [15:0] _U122_in;
wire _U122_clk;
wire [15:0] _U122_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
assign _U119_in = in[0];
assign _U119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U119 (
    .in(_U119_in),
    .clk(_U119_clk),
    .out(_U119_out)
);
assign _U120_in = in[1];
assign _U120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(_U120_in),
    .clk(_U120_clk),
    .out(_U120_out)
);
assign _U121_in = in[2];
assign _U121_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U121 (
    .in(_U121_in),
    .clk(_U121_clk),
    .out(_U121_out)
);
assign _U122_in = in[3];
assign _U122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U122 (
    .in(_U122_in),
    .clk(_U122_clk),
    .out(_U122_out)
);
assign _U123_in = in[4];
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign out[4] = _U123_out;
assign out[3] = _U122_out;
assign out[2] = _U121_out;
assign out[1] = _U120_out;
assign out[0] = _U119_out;
endmodule

module array_delay_U111 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U112_in;
wire _U112_clk;
wire [15:0] _U112_out;
wire [15:0] _U113_in;
wire _U113_clk;
wire [15:0] _U113_out;
wire [15:0] _U114_in;
wire _U114_clk;
wire [15:0] _U114_out;
wire [15:0] _U115_in;
wire _U115_clk;
wire [15:0] _U115_out;
wire [15:0] _U116_in;
wire _U116_clk;
wire [15:0] _U116_out;
assign _U112_in = in[0];
assign _U112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U112_in),
    .clk(_U112_clk),
    .out(_U112_out)
);
assign _U113_in = in[1];
assign _U113_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U113 (
    .in(_U113_in),
    .clk(_U113_clk),
    .out(_U113_out)
);
assign _U114_in = in[2];
assign _U114_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U114 (
    .in(_U114_in),
    .clk(_U114_clk),
    .out(_U114_out)
);
assign _U115_in = in[3];
assign _U115_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U115 (
    .in(_U115_in),
    .clk(_U115_clk),
    .out(_U115_out)
);
assign _U116_in = in[4];
assign _U116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U116_in),
    .clk(_U116_clk),
    .out(_U116_out)
);
assign out[4] = _U116_out;
assign out[3] = _U115_out;
assign out[2] = _U114_out;
assign out[1] = _U113_out;
assign out[0] = _U112_out;
endmodule

module array_delay_U104 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U105_in;
wire _U105_clk;
wire [15:0] _U105_out;
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire _U108_clk;
wire [15:0] _U108_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
assign _U105_in = in[0];
assign _U105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U105 (
    .in(_U105_in),
    .clk(_U105_clk),
    .out(_U105_out)
);
assign _U106_in = in[1];
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = in[2];
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = in[3];
assign _U108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U108_in),
    .clk(_U108_clk),
    .out(_U108_out)
);
assign _U109_in = in[4];
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign out[4] = _U109_out;
assign out[3] = _U108_out;
assign out[2] = _U107_out;
assign out[1] = _U106_out;
assign out[0] = _U105_out;
endmodule

module _U99_pt__U100 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U8_pt__U9 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_kernel_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
wire [15:0] _U8_in;
assign _U8_in = in0_hw_kernel_stencil[0];
_U8_pt__U9 _U8 (
    .in(_U8_in),
    .out(out_hw_kernel_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module _U83_pt__U84 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U75_pt__U76 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U6_pt__U7 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U6_in;
assign _U6_in = in0_conv_stencil[0];
_U6_pt__U7 _U6 (
    .in(_U6_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U67_pt__U68 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U612_pt__U613 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U60_pt__U61 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U598_pt__U599 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U596_pt__U597 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U593_pt__U594 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U576_pt__U577 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U573_pt__U574 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U570_pt__U571 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U568_pt__U569 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U566_pt__U567 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U550_pt__U551 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U547_pt__U548 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U543_pt__U544 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U540_pt__U541 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U53_pt__U54 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U534_pt__U535 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U531_pt__U532 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U523_pt__U524 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U520_pt__U521 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U510_pt__U511 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U507_pt__U508 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U4_pt__U5 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U4_in;
assign _U4_in = 16'h0000;
_U4_pt__U5 _U4 (
    .in(_U4_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U495_pt__U496 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U492_pt__U493 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U483_pt__U484 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U47_pt__U48 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U474_pt__U475 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U466_pt__U467 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U458_pt__U459 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U451_pt__U452 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U444_pt__U445 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U438_pt__U439 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U432_pt__U433 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U427_pt__U428 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U422_pt__U423 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U41_pt__U42 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U418_pt__U419 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U414_pt__U415 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_3_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U414_in;
wire [15:0] _U414_out;
wire [15:0] _U416_in;
wire _U416_clk;
wire [15:0] _U416_out;
wire [15:0] _U417_in;
wire _U417_clk;
wire [15:0] _U417_out;
wire [15:0] _U418_in;
wire [15:0] _U418_out;
wire [15:0] _U420_in;
wire _U420_clk;
wire [15:0] _U420_out;
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire [15:0] _U422_out;
wire [15:0] _U424_in;
wire _U424_clk;
wire [15:0] _U424_out;
wire [15:0] _U425_in;
wire _U425_clk;
wire [15:0] _U425_out;
wire [15:0] _U426_in;
wire _U426_clk;
wire [15:0] _U426_out;
wire [15:0] _U427_in;
wire [15:0] _U427_out;
wire [15:0] _U429_in;
wire _U429_clk;
wire [15:0] _U429_out;
wire [15:0] _U430_in;
wire _U430_clk;
wire [15:0] _U430_out;
wire [15:0] _U431_in;
wire _U431_clk;
wire [15:0] _U431_out;
wire [15:0] _U432_in;
wire [15:0] _U432_out;
wire [15:0] _U434_in;
wire _U434_clk;
wire [15:0] _U434_out;
wire [15:0] _U435_in;
wire _U435_clk;
wire [15:0] _U435_out;
wire [15:0] _U436_in;
wire _U436_clk;
wire [15:0] _U436_out;
wire [15:0] _U437_in;
wire _U437_clk;
wire [15:0] _U437_out;
wire [15:0] _U438_in;
wire [15:0] _U438_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire [15:0] _U444_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
wire [15:0] _U447_in;
wire _U447_clk;
wire [15:0] _U447_out;
wire [15:0] _U448_in;
wire _U448_clk;
wire [15:0] _U448_out;
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
wire [15:0] _U451_in;
wire [15:0] _U451_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
wire [15:0] _U454_in;
wire _U454_clk;
wire [15:0] _U454_out;
wire [15:0] _U455_in;
wire _U455_clk;
wire [15:0] _U455_out;
wire [15:0] _U456_in;
wire _U456_clk;
wire [15:0] _U456_out;
wire [15:0] _U457_in;
wire _U457_clk;
wire [15:0] _U457_out;
wire [15:0] _U458_in;
wire [15:0] _U458_out;
wire [15:0] _U460_in;
wire _U460_clk;
wire [15:0] _U460_out;
wire [15:0] _U461_in;
wire _U461_clk;
wire [15:0] _U461_out;
wire [15:0] _U462_in;
wire _U462_clk;
wire [15:0] _U462_out;
wire [15:0] _U463_in;
wire _U463_clk;
wire [15:0] _U463_out;
wire [15:0] _U464_in;
wire _U464_clk;
wire [15:0] _U464_out;
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire [15:0] _U466_out;
wire [15:0] _U468_in;
wire _U468_clk;
wire [15:0] _U468_out;
wire [15:0] _U469_in;
wire _U469_clk;
wire [15:0] _U469_out;
wire [15:0] _U470_in;
wire _U470_clk;
wire [15:0] _U470_out;
wire [15:0] _U471_in;
wire _U471_clk;
wire [15:0] _U471_out;
wire [15:0] _U472_in;
wire _U472_clk;
wire [15:0] _U472_out;
wire [15:0] _U473_in;
wire _U473_clk;
wire [15:0] _U473_out;
wire [15:0] _U474_in;
wire [15:0] _U474_out;
wire [15:0] _U476_in;
wire _U476_clk;
wire [15:0] _U476_out;
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire _U478_clk;
wire [15:0] _U478_out;
wire [15:0] _U479_in;
wire _U479_clk;
wire [15:0] _U479_out;
wire [15:0] _U480_in;
wire _U480_clk;
wire [15:0] _U480_out;
wire [15:0] _U481_in;
wire _U481_clk;
wire [15:0] _U481_out;
wire [15:0] _U482_in;
wire _U482_clk;
wire [15:0] _U482_out;
wire [15:0] _U483_in;
wire [15:0] _U483_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire _U487_clk;
wire [15:0] _U487_out;
wire [15:0] _U488_in;
wire _U488_clk;
wire [15:0] _U488_out;
wire [15:0] _U489_in;
wire _U489_clk;
wire [15:0] _U489_out;
wire [15:0] _U490_in;
wire _U490_clk;
wire [15:0] _U490_out;
wire [15:0] _U491_in;
wire _U491_clk;
wire [15:0] _U491_out;
wire [15:0] _U492_in;
wire [15:0] _U492_out;
wire [15:0] _U494_in;
wire _U494_clk;
wire [15:0] _U494_out;
wire [15:0] _U495_in;
wire [15:0] _U495_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
wire [15:0] _U498_in;
wire _U498_clk;
wire [15:0] _U498_out;
wire [15:0] _U499_in;
wire _U499_clk;
wire [15:0] _U499_out;
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire _U502_clk;
wire [15:0] _U502_out;
wire [15:0] _U503_in;
wire _U503_clk;
wire [15:0] _U503_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire _U506_clk;
wire [15:0] _U506_out;
wire [15:0] _U507_in;
wire [15:0] _U507_out;
wire [15:0] _U509_in;
wire _U509_clk;
wire [15:0] _U509_out;
wire [15:0] _U510_in;
wire [15:0] _U510_out;
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire _U513_clk;
wire [15:0] _U513_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
wire [15:0] _U517_in;
wire _U517_clk;
wire [15:0] _U517_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire [15:0] _U520_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire [15:0] _U523_out;
wire [15:0] _U525_in;
wire _U525_clk;
wire [15:0] _U525_out;
wire [15:0] _U526_in;
wire _U526_clk;
wire [15:0] _U526_out;
wire [15:0] _U527_in;
wire _U527_clk;
wire [15:0] _U527_out;
wire [15:0] _U528_in;
wire _U528_clk;
wire [15:0] _U528_out;
wire [15:0] _U529_in;
wire _U529_clk;
wire [15:0] _U529_out;
wire [15:0] _U530_in;
wire _U530_clk;
wire [15:0] _U530_out;
wire [15:0] _U531_in;
wire [15:0] _U531_out;
wire [15:0] _U533_in;
wire _U533_clk;
wire [15:0] _U533_out;
wire [15:0] _U534_in;
wire [15:0] _U534_out;
wire [15:0] _U536_in;
wire _U536_clk;
wire [15:0] _U536_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire _U539_clk;
wire [15:0] _U539_out;
wire [15:0] _U540_in;
wire [15:0] _U540_out;
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
wire [15:0] _U543_in;
wire [15:0] _U543_out;
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
wire [15:0] _U547_in;
wire [15:0] _U547_out;
wire [15:0] _U549_in;
wire _U549_clk;
wire [15:0] _U549_out;
wire [15:0] _U550_in;
wire [15:0] _U550_out;
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire _U553_clk;
wire [15:0] _U553_out;
wire [15:0] _U554_in;
wire _U554_clk;
wire [15:0] _U554_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
wire [15:0] _U557_in;
wire _U557_clk;
wire [15:0] _U557_out;
wire [15:0] _U558_in;
wire _U558_clk;
wire [15:0] _U558_out;
wire [15:0] _U559_in;
wire _U559_clk;
wire [15:0] _U559_out;
wire [15:0] _U560_in;
wire _U560_clk;
wire [15:0] _U560_out;
wire [15:0] _U561_in;
wire _U561_clk;
wire [15:0] _U561_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
wire [15:0] _U564_in;
wire _U564_clk;
wire [15:0] _U564_out;
wire [15:0] _U565_in;
wire _U565_clk;
wire [15:0] _U565_out;
wire [15:0] _U566_in;
wire [15:0] _U566_out;
wire [15:0] _U568_in;
wire [15:0] _U568_out;
wire [15:0] _U570_in;
wire [15:0] _U570_out;
wire [15:0] _U572_in;
wire _U572_clk;
wire [15:0] _U572_out;
wire [15:0] _U573_in;
wire [15:0] _U573_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire [15:0] _U576_out;
wire [15:0] _U578_in;
wire _U578_clk;
wire [15:0] _U578_out;
wire [15:0] _U579_in;
wire _U579_clk;
wire [15:0] _U579_out;
wire [15:0] _U580_in;
wire _U580_clk;
wire [15:0] _U580_out;
wire [15:0] _U581_in;
wire _U581_clk;
wire [15:0] _U581_out;
wire [15:0] _U582_in;
wire _U582_clk;
wire [15:0] _U582_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
wire [15:0] _U585_in;
wire _U585_clk;
wire [15:0] _U585_out;
wire [15:0] _U586_in;
wire _U586_clk;
wire [15:0] _U586_out;
wire [15:0] _U587_in;
wire _U587_clk;
wire [15:0] _U587_out;
wire [15:0] _U588_in;
wire _U588_clk;
wire [15:0] _U588_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
wire [15:0] _U592_in;
wire _U592_clk;
wire [15:0] _U592_out;
wire [15:0] _U593_in;
wire [15:0] _U593_out;
wire [15:0] _U595_in;
wire _U595_clk;
wire [15:0] _U595_out;
wire [15:0] _U596_in;
wire [15:0] _U598_in;
wire [15:0] _U598_out;
wire [15:0] _U600_in;
wire _U600_clk;
wire [15:0] _U600_out;
wire [15:0] _U601_in;
wire _U601_clk;
wire [15:0] _U601_out;
wire [15:0] _U602_in;
wire _U602_clk;
wire [15:0] _U602_out;
wire [15:0] _U603_in;
wire _U603_clk;
wire [15:0] _U603_out;
wire [15:0] _U604_in;
wire _U604_clk;
wire [15:0] _U604_out;
wire [15:0] _U605_in;
wire _U605_clk;
wire [15:0] _U605_out;
wire [15:0] _U606_in;
wire _U606_clk;
wire [15:0] _U606_out;
wire [15:0] _U607_in;
wire _U607_clk;
wire [15:0] _U607_out;
wire [15:0] _U608_in;
wire _U608_clk;
wire [15:0] _U608_out;
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
wire [15:0] _U611_in;
wire _U611_clk;
wire [15:0] _U611_out;
wire [15:0] _U612_in;
wire [15:0] _U612_out;
wire [15:0] _U614_in;
wire _U614_clk;
wire [15:0] _U614_out;
assign _U414_in = _U417_out;
_U414_pt__U415 _U414 (
    .in(_U414_in),
    .out(_U414_out)
);
assign _U416_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U416_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U416 (
    .in(_U416_in),
    .clk(_U416_clk),
    .out(_U416_out)
);
assign _U417_in = _U416_out;
assign _U417_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U417 (
    .in(_U417_in),
    .clk(_U417_clk),
    .out(_U417_out)
);
assign _U418_in = _U421_out;
_U418_pt__U419 _U418 (
    .in(_U418_in),
    .out(_U418_out)
);
assign _U420_in = in1_hw_input_global_wrapper_stencil[2];
assign _U420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U420_in),
    .clk(_U420_clk),
    .out(_U420_out)
);
assign _U421_in = _U420_out;
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = _U426_out;
_U422_pt__U423 _U422 (
    .in(_U422_in),
    .out(_U422_out)
);
assign _U424_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U424 (
    .in(_U424_in),
    .clk(_U424_clk),
    .out(_U424_out)
);
assign _U425_in = _U424_out;
assign _U425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U425 (
    .in(_U425_in),
    .clk(_U425_clk),
    .out(_U425_out)
);
assign _U426_in = _U425_out;
assign _U426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U426 (
    .in(_U426_in),
    .clk(_U426_clk),
    .out(_U426_out)
);
assign _U427_in = _U431_out;
_U427_pt__U428 _U427 (
    .in(_U427_in),
    .out(_U427_out)
);
assign _U429_in = in1_hw_input_global_wrapper_stencil[3];
assign _U429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U429 (
    .in(_U429_in),
    .clk(_U429_clk),
    .out(_U429_out)
);
assign _U430_in = _U429_out;
assign _U430_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U430 (
    .in(_U430_in),
    .clk(_U430_clk),
    .out(_U430_out)
);
assign _U431_in = _U430_out;
assign _U431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U431_in),
    .clk(_U431_clk),
    .out(_U431_out)
);
assign _U432_in = _U437_out;
_U432_pt__U433 _U432 (
    .in(_U432_in),
    .out(_U432_out)
);
assign _U434_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U434_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U434 (
    .in(_U434_in),
    .clk(_U434_clk),
    .out(_U434_out)
);
assign _U435_in = _U434_out;
assign _U435_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U435 (
    .in(_U435_in),
    .clk(_U435_clk),
    .out(_U435_out)
);
assign _U436_in = _U435_out;
assign _U436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U436 (
    .in(_U436_in),
    .clk(_U436_clk),
    .out(_U436_out)
);
assign _U437_in = _U436_out;
assign _U437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U437 (
    .in(_U437_in),
    .clk(_U437_clk),
    .out(_U437_out)
);
assign _U438_in = _U443_out;
_U438_pt__U439 _U438 (
    .in(_U438_in),
    .out(_U438_out)
);
assign _U440_in = in1_hw_input_global_wrapper_stencil[4];
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = _U440_out;
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign _U442_in = _U441_out;
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = _U442_out;
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = _U450_out;
_U444_pt__U445 _U444 (
    .in(_U444_in),
    .out(_U444_out)
);
assign _U446_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign _U447_in = _U446_out;
assign _U447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U447 (
    .in(_U447_in),
    .clk(_U447_clk),
    .out(_U447_out)
);
assign _U448_in = _U447_out;
assign _U448_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U448 (
    .in(_U448_in),
    .clk(_U448_clk),
    .out(_U448_out)
);
assign _U449_in = _U448_out;
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = _U449_out;
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign _U451_in = _U457_out;
_U451_pt__U452 _U451 (
    .in(_U451_in),
    .out(_U451_out)
);
assign _U453_in = in1_hw_input_global_wrapper_stencil[5];
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign _U454_in = _U453_out;
assign _U454_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U454 (
    .in(_U454_in),
    .clk(_U454_clk),
    .out(_U454_out)
);
assign _U455_in = _U454_out;
assign _U455_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U455 (
    .in(_U455_in),
    .clk(_U455_clk),
    .out(_U455_out)
);
assign _U456_in = _U455_out;
assign _U456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U456 (
    .in(_U456_in),
    .clk(_U456_clk),
    .out(_U456_out)
);
assign _U457_in = _U456_out;
assign _U457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U457 (
    .in(_U457_in),
    .clk(_U457_clk),
    .out(_U457_out)
);
assign _U458_in = _U465_out;
_U458_pt__U459 _U458 (
    .in(_U458_in),
    .out(_U458_out)
);
assign _U460_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U460 (
    .in(_U460_in),
    .clk(_U460_clk),
    .out(_U460_out)
);
assign _U461_in = _U460_out;
assign _U461_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U461 (
    .in(_U461_in),
    .clk(_U461_clk),
    .out(_U461_out)
);
assign _U462_in = _U461_out;
assign _U462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U462_in),
    .clk(_U462_clk),
    .out(_U462_out)
);
assign _U463_in = _U462_out;
assign _U463_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U463 (
    .in(_U463_in),
    .clk(_U463_clk),
    .out(_U463_out)
);
assign _U464_in = _U463_out;
assign _U464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U464 (
    .in(_U464_in),
    .clk(_U464_clk),
    .out(_U464_out)
);
assign _U465_in = _U464_out;
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = _U473_out;
_U466_pt__U467 _U466 (
    .in(_U466_in),
    .out(_U466_out)
);
assign _U468_in = in1_hw_input_global_wrapper_stencil[6];
assign _U468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U468_in),
    .clk(_U468_clk),
    .out(_U468_out)
);
assign _U469_in = _U468_out;
assign _U469_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U469 (
    .in(_U469_in),
    .clk(_U469_clk),
    .out(_U469_out)
);
assign _U470_in = _U469_out;
assign _U470_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U470 (
    .in(_U470_in),
    .clk(_U470_clk),
    .out(_U470_out)
);
assign _U471_in = _U470_out;
assign _U471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U471 (
    .in(_U471_in),
    .clk(_U471_clk),
    .out(_U471_out)
);
assign _U472_in = _U471_out;
assign _U472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U472 (
    .in(_U472_in),
    .clk(_U472_clk),
    .out(_U472_out)
);
assign _U473_in = _U472_out;
assign _U473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U473 (
    .in(_U473_in),
    .clk(_U473_clk),
    .out(_U473_out)
);
assign _U474_in = _U482_out;
_U474_pt__U475 _U474 (
    .in(_U474_in),
    .out(_U474_out)
);
assign _U476_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(_U476_in),
    .clk(_U476_clk),
    .out(_U476_out)
);
assign _U477_in = _U476_out;
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = _U477_out;
assign _U478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(_U478_in),
    .clk(_U478_clk),
    .out(_U478_out)
);
assign _U479_in = _U478_out;
assign _U479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(_U479_in),
    .clk(_U479_clk),
    .out(_U479_out)
);
assign _U480_in = _U479_out;
assign _U480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U480 (
    .in(_U480_in),
    .clk(_U480_clk),
    .out(_U480_out)
);
assign _U481_in = _U480_out;
assign _U481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U481_in),
    .clk(_U481_clk),
    .out(_U481_out)
);
assign _U482_in = _U481_out;
assign _U482_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U482 (
    .in(_U482_in),
    .clk(_U482_clk),
    .out(_U482_out)
);
assign _U483_in = _U491_out;
_U483_pt__U484 _U483 (
    .in(_U483_in),
    .out(_U483_out)
);
assign _U485_in = in1_hw_input_global_wrapper_stencil[7];
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = _U485_out;
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = _U486_out;
assign _U487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U487 (
    .in(_U487_in),
    .clk(_U487_clk),
    .out(_U487_out)
);
assign _U488_in = _U487_out;
assign _U488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U488 (
    .in(_U488_in),
    .clk(_U488_clk),
    .out(_U488_out)
);
assign _U489_in = _U488_out;
assign _U489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U489_in),
    .clk(_U489_clk),
    .out(_U489_out)
);
assign _U490_in = _U489_out;
assign _U490_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U490 (
    .in(_U490_in),
    .clk(_U490_clk),
    .out(_U490_out)
);
assign _U491_in = _U490_out;
assign _U491_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U491 (
    .in(_U491_in),
    .clk(_U491_clk),
    .out(_U491_out)
);
assign _U492_in = _U494_out;
_U492_pt__U493 _U492 (
    .in(_U492_in),
    .out(_U492_out)
);
assign _U494_in = 16'(_U598_out + _U612_out);
assign _U494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U494 (
    .in(_U494_in),
    .clk(_U494_clk),
    .out(_U494_out)
);
assign _U495_in = _U506_out;
_U495_pt__U496 _U495 (
    .in(_U495_in),
    .out(_U495_out)
);
assign _U497_in = 16'(_U414_out * _U418_out);
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign _U498_in = _U497_out;
assign _U498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U498_in),
    .clk(_U498_clk),
    .out(_U498_out)
);
assign _U499_in = _U498_out;
assign _U499_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(_U499_in),
    .clk(_U499_clk),
    .out(_U499_out)
);
assign _U500_in = _U499_out;
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign _U501_in = _U500_out;
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = _U501_out;
assign _U502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U502_in),
    .clk(_U502_clk),
    .out(_U502_out)
);
assign _U503_in = _U502_out;
assign _U503_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U503 (
    .in(_U503_in),
    .clk(_U503_clk),
    .out(_U503_out)
);
assign _U504_in = _U503_out;
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign _U505_in = _U504_out;
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = _U505_out;
assign _U506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U506 (
    .in(_U506_in),
    .clk(_U506_clk),
    .out(_U506_out)
);
assign _U507_in = _U509_out;
_U507_pt__U508 _U507 (
    .in(_U507_in),
    .out(_U507_out)
);
assign _U509_in = 16'(_U510_out + _U520_out);
assign _U509_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U509 (
    .in(_U509_in),
    .clk(_U509_clk),
    .out(_U509_out)
);
assign _U510_in = _U519_out;
_U510_pt__U511 _U510 (
    .in(_U510_in),
    .out(_U510_out)
);
assign _U512_in = 16'(_U422_out * _U427_out);
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = _U512_out;
assign _U513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U513_in),
    .clk(_U513_clk),
    .out(_U513_out)
);
assign _U514_in = _U513_out;
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = _U514_out;
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = _U515_out;
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign _U517_in = _U516_out;
assign _U517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(_U517_in),
    .clk(_U517_clk),
    .out(_U517_out)
);
assign _U518_in = _U517_out;
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign _U519_in = _U518_out;
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = _U522_out;
_U520_pt__U521 _U520 (
    .in(_U520_in),
    .out(_U520_out)
);
assign _U522_in = 16'(_U523_out + _U531_out);
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = _U530_out;
_U523_pt__U524 _U523 (
    .in(_U523_in),
    .out(_U523_out)
);
assign _U525_in = 16'(_U432_out * _U438_out);
assign _U525_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U525 (
    .in(_U525_in),
    .clk(_U525_clk),
    .out(_U525_out)
);
assign _U526_in = _U525_out;
assign _U526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(_U526_in),
    .clk(_U526_clk),
    .out(_U526_out)
);
assign _U527_in = _U526_out;
assign _U527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(_U527_in),
    .clk(_U527_clk),
    .out(_U527_out)
);
assign _U528_in = _U527_out;
assign _U528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(_U528_in),
    .clk(_U528_clk),
    .out(_U528_out)
);
assign _U529_in = _U528_out;
assign _U529_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U529 (
    .in(_U529_in),
    .clk(_U529_clk),
    .out(_U529_out)
);
assign _U530_in = _U529_out;
assign _U530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U530 (
    .in(_U530_in),
    .clk(_U530_clk),
    .out(_U530_out)
);
assign _U531_in = _U533_out;
_U531_pt__U532 _U531 (
    .in(_U531_in),
    .out(_U531_out)
);
assign _U533_in = 16'(_U534_out + _U540_out);
assign _U533_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U533 (
    .in(_U533_in),
    .clk(_U533_clk),
    .out(_U533_out)
);
assign _U534_in = _U539_out;
_U534_pt__U535 _U534 (
    .in(_U534_in),
    .out(_U534_out)
);
assign _U536_in = 16'(_U444_out * _U451_out);
assign _U536_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U536_in),
    .clk(_U536_clk),
    .out(_U536_out)
);
assign _U537_in = _U536_out;
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign _U538_in = _U537_out;
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = _U538_out;
assign _U539_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U539 (
    .in(_U539_in),
    .clk(_U539_clk),
    .out(_U539_out)
);
assign _U540_in = _U542_out;
_U540_pt__U541 _U540 (
    .in(_U540_in),
    .out(_U540_out)
);
assign _U542_in = 16'(_U543_out + _U547_out);
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign _U543_in = _U546_out;
_U543_pt__U544 _U543 (
    .in(_U543_in),
    .out(_U543_out)
);
assign _U545_in = 16'(_U458_out * _U466_out);
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = _U545_out;
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign _U547_in = _U549_out;
_U547_pt__U548 _U547 (
    .in(_U547_in),
    .out(_U547_out)
);
assign _U549_in = 16'(_U474_out * _U483_out);
assign _U549_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U549 (
    .in(_U549_in),
    .clk(_U549_clk),
    .out(_U549_out)
);
assign _U550_in = _U565_out;
_U550_pt__U551 _U550 (
    .in(_U550_in),
    .out(_U550_out)
);
assign _U552_in = in0_conv_stencil[0];
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = _U552_out;
assign _U553_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U553 (
    .in(_U553_in),
    .clk(_U553_clk),
    .out(_U553_out)
);
assign _U554_in = _U553_out;
assign _U554_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U554 (
    .in(_U554_in),
    .clk(_U554_clk),
    .out(_U554_out)
);
assign _U555_in = _U554_out;
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = _U555_out;
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign _U557_in = _U556_out;
assign _U557_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U557 (
    .in(_U557_in),
    .clk(_U557_clk),
    .out(_U557_out)
);
assign _U558_in = _U557_out;
assign _U558_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U558 (
    .in(_U558_in),
    .clk(_U558_clk),
    .out(_U558_out)
);
assign _U559_in = _U558_out;
assign _U559_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U559 (
    .in(_U559_in),
    .clk(_U559_clk),
    .out(_U559_out)
);
assign _U560_in = _U559_out;
assign _U560_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U560 (
    .in(_U560_in),
    .clk(_U560_clk),
    .out(_U560_out)
);
assign _U561_in = _U560_out;
assign _U561_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(_U561_in),
    .clk(_U561_clk),
    .out(_U561_out)
);
assign _U562_in = _U561_out;
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = _U562_out;
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign _U564_in = _U563_out;
assign _U564_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U564 (
    .in(_U564_in),
    .clk(_U564_clk),
    .out(_U564_out)
);
assign _U565_in = _U564_out;
assign _U565_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U565 (
    .in(_U565_in),
    .clk(_U565_clk),
    .out(_U565_out)
);
assign _U566_in = in2_hw_kernel_global_wrapper_stencil[0];
_U566_pt__U567 _U566 (
    .in(_U566_in),
    .out(_U566_out)
);
assign _U568_in = in1_hw_input_global_wrapper_stencil[0];
_U568_pt__U569 _U568 (
    .in(_U568_in),
    .out(_U568_out)
);
assign _U570_in = _U572_out;
_U570_pt__U571 _U570 (
    .in(_U570_in),
    .out(_U570_out)
);
assign _U572_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U572_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U572 (
    .in(_U572_in),
    .clk(_U572_clk),
    .out(_U572_out)
);
assign _U573_in = _U575_out;
_U573_pt__U574 _U573 (
    .in(_U573_in),
    .out(_U573_out)
);
assign _U575_in = in1_hw_input_global_wrapper_stencil[1];
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = _U592_out;
_U576_pt__U577 _U576 (
    .in(_U576_in),
    .out(_U576_out)
);
assign _U578_in = 16'(_U566_out * _U568_out);
assign _U578_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U578 (
    .in(_U578_in),
    .clk(_U578_clk),
    .out(_U578_out)
);
assign _U579_in = _U578_out;
assign _U579_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U579 (
    .in(_U579_in),
    .clk(_U579_clk),
    .out(_U579_out)
);
assign _U580_in = _U579_out;
assign _U580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U580_in),
    .clk(_U580_clk),
    .out(_U580_out)
);
assign _U581_in = _U580_out;
assign _U581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U581_in),
    .clk(_U581_clk),
    .out(_U581_out)
);
assign _U582_in = _U581_out;
assign _U582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U582_in),
    .clk(_U582_clk),
    .out(_U582_out)
);
assign _U583_in = _U582_out;
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = _U583_out;
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign _U585_in = _U584_out;
assign _U585_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U585 (
    .in(_U585_in),
    .clk(_U585_clk),
    .out(_U585_out)
);
assign _U586_in = _U585_out;
assign _U586_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U586 (
    .in(_U586_in),
    .clk(_U586_clk),
    .out(_U586_out)
);
assign _U587_in = _U586_out;
assign _U587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U587_in),
    .clk(_U587_clk),
    .out(_U587_out)
);
assign _U588_in = _U587_out;
assign _U588_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U588 (
    .in(_U588_in),
    .clk(_U588_clk),
    .out(_U588_out)
);
assign _U589_in = _U588_out;
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = _U589_out;
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = _U590_out;
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign _U592_in = _U591_out;
assign _U592_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U592 (
    .in(_U592_in),
    .clk(_U592_clk),
    .out(_U592_out)
);
assign _U593_in = _U595_out;
_U593_pt__U594 _U593 (
    .in(_U593_in),
    .out(_U593_out)
);
assign _U595_in = 16'(_U550_out + _U492_out);
assign _U595_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U595 (
    .in(_U595_in),
    .clk(_U595_clk),
    .out(_U595_out)
);
assign _U596_in = 16'(_U576_out + _U593_out);
_U596_pt__U597 _U596 (
    .in(_U596_in),
    .out(out_conv_stencil)
);
assign _U598_in = _U611_out;
_U598_pt__U599 _U598 (
    .in(_U598_in),
    .out(_U598_out)
);
assign _U600_in = 16'(_U570_out * _U573_out);
assign _U600_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U600 (
    .in(_U600_in),
    .clk(_U600_clk),
    .out(_U600_out)
);
assign _U601_in = _U600_out;
assign _U601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U601_in),
    .clk(_U601_clk),
    .out(_U601_out)
);
assign _U602_in = _U601_out;
assign _U602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U602_in),
    .clk(_U602_clk),
    .out(_U602_out)
);
assign _U603_in = _U602_out;
assign _U603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U603 (
    .in(_U603_in),
    .clk(_U603_clk),
    .out(_U603_out)
);
assign _U604_in = _U603_out;
assign _U604_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U604 (
    .in(_U604_in),
    .clk(_U604_clk),
    .out(_U604_out)
);
assign _U605_in = _U604_out;
assign _U605_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U605 (
    .in(_U605_in),
    .clk(_U605_clk),
    .out(_U605_out)
);
assign _U606_in = _U605_out;
assign _U606_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U606 (
    .in(_U606_in),
    .clk(_U606_clk),
    .out(_U606_out)
);
assign _U607_in = _U606_out;
assign _U607_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U607 (
    .in(_U607_in),
    .clk(_U607_clk),
    .out(_U607_out)
);
assign _U608_in = _U607_out;
assign _U608_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U608 (
    .in(_U608_in),
    .clk(_U608_clk),
    .out(_U608_out)
);
assign _U609_in = _U608_out;
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = _U609_out;
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
assign _U611_in = _U610_out;
assign _U611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U611 (
    .in(_U611_in),
    .clk(_U611_clk),
    .out(_U611_out)
);
assign _U612_in = _U614_out;
_U612_pt__U613 _U612 (
    .in(_U612_in),
    .out(_U612_out)
);
assign _U614_in = 16'(_U495_out + _U507_out);
assign _U614_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U614 (
    .in(_U614_in),
    .clk(_U614_clk),
    .out(_U614_out)
);
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U412_pt__U413 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_2_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U412_in;
assign _U412_in = 16'h0000;
_U412_pt__U413 _U412 (
    .in(_U412_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U404_pt__U405 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U396_pt__U397 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U389_pt__U390 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U382_pt__U383 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U376_pt__U377 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U370_pt__U371 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U36_pt__U37 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U365_pt__U366 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U360_pt__U361 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U356_pt__U357 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U352_pt__U353 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U349_pt__U350 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U346_pt__U347 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U344_pt__U345 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U342_pt__U343 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U326_pt__U327 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U31_pt__U32 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U310_pt__U311 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U2_pt__U3 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_1_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U2_in;
assign _U2_in = 16'h0000;
_U2_pt__U3 _U2 (
    .in(_U2_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U295_pt__U296 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U292_pt__U293 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U288_pt__U289 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U285_pt__U286 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U27_pt__U28 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U279_pt__U280 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U276_pt__U277 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U268_pt__U269 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U265_pt__U266 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U255_pt__U256 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U252_pt__U253 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U240_pt__U241 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U23_pt__U24 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U237_pt__U238 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U234_pt__U235 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U220_pt__U221 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U218_pt__U219 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U214_pt__U215 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U211_pt__U212 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_5_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U211_in;
wire [15:0] _U211_out;
wire [15:0] _U213_in;
wire _U213_clk;
wire [15:0] _U213_out;
wire [15:0] _U214_in;
wire [15:0] _U214_out;
wire [15:0] _U216_in;
wire _U216_clk;
wire [15:0] _U216_out;
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire [15:0] _U220_in;
wire [15:0] _U220_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
wire [15:0] _U223_in;
wire _U223_clk;
wire [15:0] _U223_out;
wire [15:0] _U224_in;
wire _U224_clk;
wire [15:0] _U224_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
wire [15:0] _U229_in;
wire _U229_clk;
wire [15:0] _U229_out;
wire [15:0] _U230_in;
wire _U230_clk;
wire [15:0] _U230_out;
wire [15:0] _U231_in;
wire _U231_clk;
wire [15:0] _U231_out;
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
wire [15:0] _U233_in;
wire _U233_clk;
wire [15:0] _U233_out;
wire [15:0] _U234_in;
wire [15:0] _U234_out;
wire [15:0] _U236_in;
wire _U236_clk;
wire [15:0] _U236_out;
wire [15:0] _U237_in;
wire [15:0] _U237_out;
wire [15:0] _U239_in;
wire _U239_clk;
wire [15:0] _U239_out;
wire [15:0] _U240_in;
wire [15:0] _U240_out;
wire [15:0] _U242_in;
wire _U242_clk;
wire [15:0] _U242_out;
wire [15:0] _U243_in;
wire _U243_clk;
wire [15:0] _U243_out;
wire [15:0] _U244_in;
wire _U244_clk;
wire [15:0] _U244_out;
wire [15:0] _U245_in;
wire _U245_clk;
wire [15:0] _U245_out;
wire [15:0] _U246_in;
wire _U246_clk;
wire [15:0] _U246_out;
wire [15:0] _U247_in;
wire _U247_clk;
wire [15:0] _U247_out;
wire [15:0] _U248_in;
wire _U248_clk;
wire [15:0] _U248_out;
wire [15:0] _U249_in;
wire _U249_clk;
wire [15:0] _U249_out;
wire [15:0] _U250_in;
wire _U250_clk;
wire [15:0] _U250_out;
wire [15:0] _U251_in;
wire _U251_clk;
wire [15:0] _U251_out;
wire [15:0] _U252_in;
wire [15:0] _U252_out;
wire [15:0] _U254_in;
wire _U254_clk;
wire [15:0] _U254_out;
wire [15:0] _U255_in;
wire [15:0] _U255_out;
wire [15:0] _U257_in;
wire _U257_clk;
wire [15:0] _U257_out;
wire [15:0] _U258_in;
wire _U258_clk;
wire [15:0] _U258_out;
wire [15:0] _U259_in;
wire _U259_clk;
wire [15:0] _U259_out;
wire [15:0] _U260_in;
wire _U260_clk;
wire [15:0] _U260_out;
wire [15:0] _U261_in;
wire _U261_clk;
wire [15:0] _U261_out;
wire [15:0] _U262_in;
wire _U262_clk;
wire [15:0] _U262_out;
wire [15:0] _U263_in;
wire _U263_clk;
wire [15:0] _U263_out;
wire [15:0] _U264_in;
wire _U264_clk;
wire [15:0] _U264_out;
wire [15:0] _U265_in;
wire [15:0] _U265_out;
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire [15:0] _U268_out;
wire [15:0] _U270_in;
wire _U270_clk;
wire [15:0] _U270_out;
wire [15:0] _U271_in;
wire _U271_clk;
wire [15:0] _U271_out;
wire [15:0] _U272_in;
wire _U272_clk;
wire [15:0] _U272_out;
wire [15:0] _U273_in;
wire _U273_clk;
wire [15:0] _U273_out;
wire [15:0] _U274_in;
wire _U274_clk;
wire [15:0] _U274_out;
wire [15:0] _U275_in;
wire _U275_clk;
wire [15:0] _U275_out;
wire [15:0] _U276_in;
wire [15:0] _U276_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire [15:0] _U279_out;
wire [15:0] _U281_in;
wire _U281_clk;
wire [15:0] _U281_out;
wire [15:0] _U282_in;
wire _U282_clk;
wire [15:0] _U282_out;
wire [15:0] _U283_in;
wire _U283_clk;
wire [15:0] _U283_out;
wire [15:0] _U284_in;
wire _U284_clk;
wire [15:0] _U284_out;
wire [15:0] _U285_in;
wire [15:0] _U285_out;
wire [15:0] _U287_in;
wire _U287_clk;
wire [15:0] _U287_out;
wire [15:0] _U288_in;
wire [15:0] _U288_out;
wire [15:0] _U290_in;
wire _U290_clk;
wire [15:0] _U290_out;
wire [15:0] _U291_in;
wire _U291_clk;
wire [15:0] _U291_out;
wire [15:0] _U292_in;
wire [15:0] _U292_out;
wire [15:0] _U294_in;
wire _U294_clk;
wire [15:0] _U294_out;
wire [15:0] _U295_in;
wire [15:0] _U295_out;
wire [15:0] _U297_in;
wire _U297_clk;
wire [15:0] _U297_out;
wire [15:0] _U298_in;
wire _U298_clk;
wire [15:0] _U298_out;
wire [15:0] _U299_in;
wire _U299_clk;
wire [15:0] _U299_out;
wire [15:0] _U300_in;
wire _U300_clk;
wire [15:0] _U300_out;
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire _U303_clk;
wire [15:0] _U303_out;
wire [15:0] _U304_in;
wire _U304_clk;
wire [15:0] _U304_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
wire [15:0] _U306_in;
wire _U306_clk;
wire [15:0] _U306_out;
wire [15:0] _U307_in;
wire _U307_clk;
wire [15:0] _U307_out;
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire [15:0] _U310_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
wire [15:0] _U313_in;
wire _U313_clk;
wire [15:0] _U313_out;
wire [15:0] _U314_in;
wire _U314_clk;
wire [15:0] _U314_out;
wire [15:0] _U315_in;
wire _U315_clk;
wire [15:0] _U315_out;
wire [15:0] _U316_in;
wire _U316_clk;
wire [15:0] _U316_out;
wire [15:0] _U317_in;
wire _U317_clk;
wire [15:0] _U317_out;
wire [15:0] _U318_in;
wire _U318_clk;
wire [15:0] _U318_out;
wire [15:0] _U319_in;
wire _U319_clk;
wire [15:0] _U319_out;
wire [15:0] _U320_in;
wire _U320_clk;
wire [15:0] _U320_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire _U322_clk;
wire [15:0] _U322_out;
wire [15:0] _U323_in;
wire _U323_clk;
wire [15:0] _U323_out;
wire [15:0] _U324_in;
wire _U324_clk;
wire [15:0] _U324_out;
wire [15:0] _U325_in;
wire _U325_clk;
wire [15:0] _U325_out;
wire [15:0] _U326_in;
wire [15:0] _U326_out;
wire [15:0] _U328_in;
wire _U328_clk;
wire [15:0] _U328_out;
wire [15:0] _U329_in;
wire _U329_clk;
wire [15:0] _U329_out;
wire [15:0] _U330_in;
wire _U330_clk;
wire [15:0] _U330_out;
wire [15:0] _U331_in;
wire _U331_clk;
wire [15:0] _U331_out;
wire [15:0] _U332_in;
wire _U332_clk;
wire [15:0] _U332_out;
wire [15:0] _U333_in;
wire _U333_clk;
wire [15:0] _U333_out;
wire [15:0] _U334_in;
wire _U334_clk;
wire [15:0] _U334_out;
wire [15:0] _U335_in;
wire _U335_clk;
wire [15:0] _U335_out;
wire [15:0] _U336_in;
wire _U336_clk;
wire [15:0] _U336_out;
wire [15:0] _U337_in;
wire _U337_clk;
wire [15:0] _U337_out;
wire [15:0] _U338_in;
wire _U338_clk;
wire [15:0] _U338_out;
wire [15:0] _U339_in;
wire _U339_clk;
wire [15:0] _U339_out;
wire [15:0] _U340_in;
wire _U340_clk;
wire [15:0] _U340_out;
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire [15:0] _U342_out;
wire [15:0] _U344_in;
wire [15:0] _U344_out;
wire [15:0] _U346_in;
wire [15:0] _U346_out;
wire [15:0] _U348_in;
wire _U348_clk;
wire [15:0] _U348_out;
wire [15:0] _U349_in;
wire [15:0] _U349_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire [15:0] _U352_out;
wire [15:0] _U354_in;
wire _U354_clk;
wire [15:0] _U354_out;
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire [15:0] _U356_out;
wire [15:0] _U358_in;
wire _U358_clk;
wire [15:0] _U358_out;
wire [15:0] _U359_in;
wire _U359_clk;
wire [15:0] _U359_out;
wire [15:0] _U360_in;
wire [15:0] _U360_out;
wire [15:0] _U362_in;
wire _U362_clk;
wire [15:0] _U362_out;
wire [15:0] _U363_in;
wire _U363_clk;
wire [15:0] _U363_out;
wire [15:0] _U364_in;
wire _U364_clk;
wire [15:0] _U364_out;
wire [15:0] _U365_in;
wire [15:0] _U365_out;
wire [15:0] _U367_in;
wire _U367_clk;
wire [15:0] _U367_out;
wire [15:0] _U368_in;
wire _U368_clk;
wire [15:0] _U368_out;
wire [15:0] _U369_in;
wire _U369_clk;
wire [15:0] _U369_out;
wire [15:0] _U370_in;
wire [15:0] _U370_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire _U373_clk;
wire [15:0] _U373_out;
wire [15:0] _U374_in;
wire _U374_clk;
wire [15:0] _U374_out;
wire [15:0] _U375_in;
wire _U375_clk;
wire [15:0] _U375_out;
wire [15:0] _U376_in;
wire [15:0] _U376_out;
wire [15:0] _U378_in;
wire _U378_clk;
wire [15:0] _U378_out;
wire [15:0] _U379_in;
wire _U379_clk;
wire [15:0] _U379_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
wire [15:0] _U381_in;
wire _U381_clk;
wire [15:0] _U381_out;
wire [15:0] _U382_in;
wire [15:0] _U382_out;
wire [15:0] _U384_in;
wire _U384_clk;
wire [15:0] _U384_out;
wire [15:0] _U385_in;
wire _U385_clk;
wire [15:0] _U385_out;
wire [15:0] _U386_in;
wire _U386_clk;
wire [15:0] _U386_out;
wire [15:0] _U387_in;
wire _U387_clk;
wire [15:0] _U387_out;
wire [15:0] _U388_in;
wire _U388_clk;
wire [15:0] _U388_out;
wire [15:0] _U389_in;
wire [15:0] _U389_out;
wire [15:0] _U391_in;
wire _U391_clk;
wire [15:0] _U391_out;
wire [15:0] _U392_in;
wire _U392_clk;
wire [15:0] _U392_out;
wire [15:0] _U393_in;
wire _U393_clk;
wire [15:0] _U393_out;
wire [15:0] _U394_in;
wire _U394_clk;
wire [15:0] _U394_out;
wire [15:0] _U395_in;
wire _U395_clk;
wire [15:0] _U395_out;
wire [15:0] _U396_in;
wire [15:0] _U396_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
wire [15:0] _U400_in;
wire _U400_clk;
wire [15:0] _U400_out;
wire [15:0] _U401_in;
wire _U401_clk;
wire [15:0] _U401_out;
wire [15:0] _U402_in;
wire _U402_clk;
wire [15:0] _U402_out;
wire [15:0] _U403_in;
wire _U403_clk;
wire [15:0] _U403_out;
wire [15:0] _U404_in;
wire [15:0] _U404_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire _U407_clk;
wire [15:0] _U407_out;
wire [15:0] _U408_in;
wire _U408_clk;
wire [15:0] _U408_out;
wire [15:0] _U409_in;
wire _U409_clk;
wire [15:0] _U409_out;
wire [15:0] _U410_in;
wire _U410_clk;
wire [15:0] _U410_out;
wire [15:0] _U411_in;
wire _U411_clk;
wire [15:0] _U411_out;
assign _U211_in = _U213_out;
_U211_pt__U212 _U211 (
    .in(_U211_in),
    .out(_U211_out)
);
assign _U213_in = 16'(_U310_out * _U326_out);
assign _U213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(_U213_in),
    .clk(_U213_clk),
    .out(_U213_out)
);
assign _U214_in = _U217_out;
_U214_pt__U215 _U214 (
    .in(_U214_in),
    .out(_U214_out)
);
assign _U216_in = 16'(_U295_out + _U237_out);
assign _U216_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(_U216_in),
    .clk(_U216_clk),
    .out(_U216_out)
);
assign _U217_in = _U216_out;
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = 16'(_U211_out + _U214_out);
_U218_pt__U219 _U218 (
    .in(_U218_in),
    .out(out_conv_stencil)
);
assign _U220_in = _U233_out;
_U220_pt__U221 _U220 (
    .in(_U220_in),
    .out(_U220_out)
);
assign _U222_in = 16'(_U342_out * _U344_out);
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign _U223_in = _U222_out;
assign _U223_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U223 (
    .in(_U223_in),
    .clk(_U223_clk),
    .out(_U223_out)
);
assign _U224_in = _U223_out;
assign _U224_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U224 (
    .in(_U224_in),
    .clk(_U224_clk),
    .out(_U224_out)
);
assign _U225_in = _U224_out;
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = _U225_out;
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = _U226_out;
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = _U227_out;
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign _U229_in = _U228_out;
assign _U229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U229_in),
    .clk(_U229_clk),
    .out(_U229_out)
);
assign _U230_in = _U229_out;
assign _U230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U230 (
    .in(_U230_in),
    .clk(_U230_clk),
    .out(_U230_out)
);
assign _U231_in = _U230_out;
assign _U231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U231 (
    .in(_U231_in),
    .clk(_U231_clk),
    .out(_U231_out)
);
assign _U232_in = _U231_out;
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign _U233_in = _U232_out;
assign _U233_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U233 (
    .in(_U233_in),
    .clk(_U233_clk),
    .out(_U233_out)
);
assign _U234_in = _U236_out;
_U234_pt__U235 _U234 (
    .in(_U234_in),
    .out(_U234_out)
);
assign _U236_in = 16'(_U240_out + _U252_out);
assign _U236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U236 (
    .in(_U236_in),
    .clk(_U236_clk),
    .out(_U236_out)
);
assign _U237_in = _U239_out;
_U237_pt__U238 _U237 (
    .in(_U237_in),
    .out(_U237_out)
);
assign _U239_in = 16'(_U220_out + _U234_out);
assign _U239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U239 (
    .in(_U239_in),
    .clk(_U239_clk),
    .out(_U239_out)
);
assign _U240_in = _U251_out;
_U240_pt__U241 _U240 (
    .in(_U240_in),
    .out(_U240_out)
);
assign _U242_in = 16'(_U346_out * _U349_out);
assign _U242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U242_in),
    .clk(_U242_clk),
    .out(_U242_out)
);
assign _U243_in = _U242_out;
assign _U243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U243_in),
    .clk(_U243_clk),
    .out(_U243_out)
);
assign _U244_in = _U243_out;
assign _U244_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U244 (
    .in(_U244_in),
    .clk(_U244_clk),
    .out(_U244_out)
);
assign _U245_in = _U244_out;
assign _U245_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U245 (
    .in(_U245_in),
    .clk(_U245_clk),
    .out(_U245_out)
);
assign _U246_in = _U245_out;
assign _U246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(_U246_in),
    .clk(_U246_clk),
    .out(_U246_out)
);
assign _U247_in = _U246_out;
assign _U247_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U247 (
    .in(_U247_in),
    .clk(_U247_clk),
    .out(_U247_out)
);
assign _U248_in = _U247_out;
assign _U248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U248 (
    .in(_U248_in),
    .clk(_U248_clk),
    .out(_U248_out)
);
assign _U249_in = _U248_out;
assign _U249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U249 (
    .in(_U249_in),
    .clk(_U249_clk),
    .out(_U249_out)
);
assign _U250_in = _U249_out;
assign _U250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U250 (
    .in(_U250_in),
    .clk(_U250_clk),
    .out(_U250_out)
);
assign _U251_in = _U250_out;
assign _U251_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U251 (
    .in(_U251_in),
    .clk(_U251_clk),
    .out(_U251_out)
);
assign _U252_in = _U254_out;
_U252_pt__U253 _U252 (
    .in(_U252_in),
    .out(_U252_out)
);
assign _U254_in = 16'(_U255_out + _U265_out);
assign _U254_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U254 (
    .in(_U254_in),
    .clk(_U254_clk),
    .out(_U254_out)
);
assign _U255_in = _U264_out;
_U255_pt__U256 _U255 (
    .in(_U255_in),
    .out(_U255_out)
);
assign _U257_in = 16'(_U352_out * _U356_out);
assign _U257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U257 (
    .in(_U257_in),
    .clk(_U257_clk),
    .out(_U257_out)
);
assign _U258_in = _U257_out;
assign _U258_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U258 (
    .in(_U258_in),
    .clk(_U258_clk),
    .out(_U258_out)
);
assign _U259_in = _U258_out;
assign _U259_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U259 (
    .in(_U259_in),
    .clk(_U259_clk),
    .out(_U259_out)
);
assign _U260_in = _U259_out;
assign _U260_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U260_in),
    .clk(_U260_clk),
    .out(_U260_out)
);
assign _U261_in = _U260_out;
assign _U261_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U261 (
    .in(_U261_in),
    .clk(_U261_clk),
    .out(_U261_out)
);
assign _U262_in = _U261_out;
assign _U262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U262 (
    .in(_U262_in),
    .clk(_U262_clk),
    .out(_U262_out)
);
assign _U263_in = _U262_out;
assign _U263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U263 (
    .in(_U263_in),
    .clk(_U263_clk),
    .out(_U263_out)
);
assign _U264_in = _U263_out;
assign _U264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U264_in),
    .clk(_U264_clk),
    .out(_U264_out)
);
assign _U265_in = _U267_out;
_U265_pt__U266 _U265 (
    .in(_U265_in),
    .out(_U265_out)
);
assign _U267_in = 16'(_U268_out + _U276_out);
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = _U275_out;
_U268_pt__U269 _U268 (
    .in(_U268_in),
    .out(_U268_out)
);
assign _U270_in = 16'(_U360_out * _U365_out);
assign _U270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(_U270_in),
    .clk(_U270_clk),
    .out(_U270_out)
);
assign _U271_in = _U270_out;
assign _U271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U271_in),
    .clk(_U271_clk),
    .out(_U271_out)
);
assign _U272_in = _U271_out;
assign _U272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U272_in),
    .clk(_U272_clk),
    .out(_U272_out)
);
assign _U273_in = _U272_out;
assign _U273_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U273 (
    .in(_U273_in),
    .clk(_U273_clk),
    .out(_U273_out)
);
assign _U274_in = _U273_out;
assign _U274_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U274 (
    .in(_U274_in),
    .clk(_U274_clk),
    .out(_U274_out)
);
assign _U275_in = _U274_out;
assign _U275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U275 (
    .in(_U275_in),
    .clk(_U275_clk),
    .out(_U275_out)
);
assign _U276_in = _U278_out;
_U276_pt__U277 _U276 (
    .in(_U276_in),
    .out(_U276_out)
);
assign _U278_in = 16'(_U279_out + _U285_out);
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = _U284_out;
_U279_pt__U280 _U279 (
    .in(_U279_in),
    .out(_U279_out)
);
assign _U281_in = 16'(_U370_out * _U376_out);
assign _U281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U281_in),
    .clk(_U281_clk),
    .out(_U281_out)
);
assign _U282_in = _U281_out;
assign _U282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U282 (
    .in(_U282_in),
    .clk(_U282_clk),
    .out(_U282_out)
);
assign _U283_in = _U282_out;
assign _U283_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U283 (
    .in(_U283_in),
    .clk(_U283_clk),
    .out(_U283_out)
);
assign _U284_in = _U283_out;
assign _U284_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U284 (
    .in(_U284_in),
    .clk(_U284_clk),
    .out(_U284_out)
);
assign _U285_in = _U287_out;
_U285_pt__U286 _U285 (
    .in(_U285_in),
    .out(_U285_out)
);
assign _U287_in = 16'(_U288_out + _U292_out);
assign _U287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U287 (
    .in(_U287_in),
    .clk(_U287_clk),
    .out(_U287_out)
);
assign _U288_in = _U291_out;
_U288_pt__U289 _U288 (
    .in(_U288_in),
    .out(_U288_out)
);
assign _U290_in = 16'(_U382_out * _U389_out);
assign _U290_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U290 (
    .in(_U290_in),
    .clk(_U290_clk),
    .out(_U290_out)
);
assign _U291_in = _U290_out;
assign _U291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U291 (
    .in(_U291_in),
    .clk(_U291_clk),
    .out(_U291_out)
);
assign _U292_in = _U294_out;
_U292_pt__U293 _U292 (
    .in(_U292_in),
    .out(_U292_out)
);
assign _U294_in = 16'(_U396_out * _U404_out);
assign _U294_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U294 (
    .in(_U294_in),
    .clk(_U294_clk),
    .out(_U294_out)
);
assign _U295_in = _U309_out;
_U295_pt__U296 _U295 (
    .in(_U295_in),
    .out(_U295_out)
);
assign _U297_in = in0_conv_stencil[0];
assign _U297_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U297 (
    .in(_U297_in),
    .clk(_U297_clk),
    .out(_U297_out)
);
assign _U298_in = _U297_out;
assign _U298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U298 (
    .in(_U298_in),
    .clk(_U298_clk),
    .out(_U298_out)
);
assign _U299_in = _U298_out;
assign _U299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U299_in),
    .clk(_U299_clk),
    .out(_U299_out)
);
assign _U300_in = _U299_out;
assign _U300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U300 (
    .in(_U300_in),
    .clk(_U300_clk),
    .out(_U300_out)
);
assign _U301_in = _U300_out;
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = _U301_out;
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = _U302_out;
assign _U303_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U303 (
    .in(_U303_in),
    .clk(_U303_clk),
    .out(_U303_out)
);
assign _U304_in = _U303_out;
assign _U304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U304 (
    .in(_U304_in),
    .clk(_U304_clk),
    .out(_U304_out)
);
assign _U305_in = _U304_out;
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign _U306_in = _U305_out;
assign _U306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U306_in),
    .clk(_U306_clk),
    .out(_U306_out)
);
assign _U307_in = _U306_out;
assign _U307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U307 (
    .in(_U307_in),
    .clk(_U307_clk),
    .out(_U307_out)
);
assign _U308_in = _U307_out;
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = _U308_out;
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = _U325_out;
_U310_pt__U311 _U310 (
    .in(_U310_in),
    .out(_U310_out)
);
assign _U312_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign _U313_in = _U312_out;
assign _U313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U313 (
    .in(_U313_in),
    .clk(_U313_clk),
    .out(_U313_out)
);
assign _U314_in = _U313_out;
assign _U314_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U314 (
    .in(_U314_in),
    .clk(_U314_clk),
    .out(_U314_out)
);
assign _U315_in = _U314_out;
assign _U315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U315_in),
    .clk(_U315_clk),
    .out(_U315_out)
);
assign _U316_in = _U315_out;
assign _U316_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U316 (
    .in(_U316_in),
    .clk(_U316_clk),
    .out(_U316_out)
);
assign _U317_in = _U316_out;
assign _U317_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U317 (
    .in(_U317_in),
    .clk(_U317_clk),
    .out(_U317_out)
);
assign _U318_in = _U317_out;
assign _U318_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U318 (
    .in(_U318_in),
    .clk(_U318_clk),
    .out(_U318_out)
);
assign _U319_in = _U318_out;
assign _U319_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U319 (
    .in(_U319_in),
    .clk(_U319_clk),
    .out(_U319_out)
);
assign _U320_in = _U319_out;
assign _U320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U320_in),
    .clk(_U320_clk),
    .out(_U320_out)
);
assign _U321_in = _U320_out;
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = _U321_out;
assign _U322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U322 (
    .in(_U322_in),
    .clk(_U322_clk),
    .out(_U322_out)
);
assign _U323_in = _U322_out;
assign _U323_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U323 (
    .in(_U323_in),
    .clk(_U323_clk),
    .out(_U323_out)
);
assign _U324_in = _U323_out;
assign _U324_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U324 (
    .in(_U324_in),
    .clk(_U324_clk),
    .out(_U324_out)
);
assign _U325_in = _U324_out;
assign _U325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U325 (
    .in(_U325_in),
    .clk(_U325_clk),
    .out(_U325_out)
);
assign _U326_in = _U341_out;
_U326_pt__U327 _U326 (
    .in(_U326_in),
    .out(_U326_out)
);
assign _U328_in = in1_hw_input_global_wrapper_stencil[0];
assign _U328_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U328 (
    .in(_U328_in),
    .clk(_U328_clk),
    .out(_U328_out)
);
assign _U329_in = _U328_out;
assign _U329_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U329 (
    .in(_U329_in),
    .clk(_U329_clk),
    .out(_U329_out)
);
assign _U330_in = _U329_out;
assign _U330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U330_in),
    .clk(_U330_clk),
    .out(_U330_out)
);
assign _U331_in = _U330_out;
assign _U331_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U331 (
    .in(_U331_in),
    .clk(_U331_clk),
    .out(_U331_out)
);
assign _U332_in = _U331_out;
assign _U332_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U332 (
    .in(_U332_in),
    .clk(_U332_clk),
    .out(_U332_out)
);
assign _U333_in = _U332_out;
assign _U333_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U333 (
    .in(_U333_in),
    .clk(_U333_clk),
    .out(_U333_out)
);
assign _U334_in = _U333_out;
assign _U334_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U334 (
    .in(_U334_in),
    .clk(_U334_clk),
    .out(_U334_out)
);
assign _U335_in = _U334_out;
assign _U335_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U335 (
    .in(_U335_in),
    .clk(_U335_clk),
    .out(_U335_out)
);
assign _U336_in = _U335_out;
assign _U336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(_U336_in),
    .clk(_U336_clk),
    .out(_U336_out)
);
assign _U337_in = _U336_out;
assign _U337_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U337 (
    .in(_U337_in),
    .clk(_U337_clk),
    .out(_U337_out)
);
assign _U338_in = _U337_out;
assign _U338_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U338 (
    .in(_U338_in),
    .clk(_U338_clk),
    .out(_U338_out)
);
assign _U339_in = _U338_out;
assign _U339_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U339 (
    .in(_U339_in),
    .clk(_U339_clk),
    .out(_U339_out)
);
assign _U340_in = _U339_out;
assign _U340_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U340 (
    .in(_U340_in),
    .clk(_U340_clk),
    .out(_U340_out)
);
assign _U341_in = _U340_out;
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = in2_hw_kernel_global_wrapper_stencil[1];
_U342_pt__U343 _U342 (
    .in(_U342_in),
    .out(_U342_out)
);
assign _U344_in = in1_hw_input_global_wrapper_stencil[1];
_U344_pt__U345 _U344 (
    .in(_U344_in),
    .out(_U344_out)
);
assign _U346_in = _U348_out;
_U346_pt__U347 _U346 (
    .in(_U346_in),
    .out(_U346_out)
);
assign _U348_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U348_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U348 (
    .in(_U348_in),
    .clk(_U348_clk),
    .out(_U348_out)
);
assign _U349_in = _U351_out;
_U349_pt__U350 _U349 (
    .in(_U349_in),
    .out(_U349_out)
);
assign _U351_in = in1_hw_input_global_wrapper_stencil[2];
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = _U355_out;
_U352_pt__U353 _U352 (
    .in(_U352_in),
    .out(_U352_out)
);
assign _U354_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U354_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U354 (
    .in(_U354_in),
    .clk(_U354_clk),
    .out(_U354_out)
);
assign _U355_in = _U354_out;
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = _U359_out;
_U356_pt__U357 _U356 (
    .in(_U356_in),
    .out(_U356_out)
);
assign _U358_in = in1_hw_input_global_wrapper_stencil[3];
assign _U358_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U358 (
    .in(_U358_in),
    .clk(_U358_clk),
    .out(_U358_out)
);
assign _U359_in = _U358_out;
assign _U359_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U359 (
    .in(_U359_in),
    .clk(_U359_clk),
    .out(_U359_out)
);
assign _U360_in = _U364_out;
_U360_pt__U361 _U360 (
    .in(_U360_in),
    .out(_U360_out)
);
assign _U362_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U362_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U362 (
    .in(_U362_in),
    .clk(_U362_clk),
    .out(_U362_out)
);
assign _U363_in = _U362_out;
assign _U363_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U363 (
    .in(_U363_in),
    .clk(_U363_clk),
    .out(_U363_out)
);
assign _U364_in = _U363_out;
assign _U364_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U364 (
    .in(_U364_in),
    .clk(_U364_clk),
    .out(_U364_out)
);
assign _U365_in = _U369_out;
_U365_pt__U366 _U365 (
    .in(_U365_in),
    .out(_U365_out)
);
assign _U367_in = in1_hw_input_global_wrapper_stencil[4];
assign _U367_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U367 (
    .in(_U367_in),
    .clk(_U367_clk),
    .out(_U367_out)
);
assign _U368_in = _U367_out;
assign _U368_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U368 (
    .in(_U368_in),
    .clk(_U368_clk),
    .out(_U368_out)
);
assign _U369_in = _U368_out;
assign _U369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U369 (
    .in(_U369_in),
    .clk(_U369_clk),
    .out(_U369_out)
);
assign _U370_in = _U375_out;
_U370_pt__U371 _U370 (
    .in(_U370_in),
    .out(_U370_out)
);
assign _U372_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = _U372_out;
assign _U373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U373 (
    .in(_U373_in),
    .clk(_U373_clk),
    .out(_U373_out)
);
assign _U374_in = _U373_out;
assign _U374_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U374 (
    .in(_U374_in),
    .clk(_U374_clk),
    .out(_U374_out)
);
assign _U375_in = _U374_out;
assign _U375_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U375 (
    .in(_U375_in),
    .clk(_U375_clk),
    .out(_U375_out)
);
assign _U376_in = _U381_out;
_U376_pt__U377 _U376 (
    .in(_U376_in),
    .out(_U376_out)
);
assign _U378_in = in1_hw_input_global_wrapper_stencil[5];
assign _U378_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U378 (
    .in(_U378_in),
    .clk(_U378_clk),
    .out(_U378_out)
);
assign _U379_in = _U378_out;
assign _U379_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U379 (
    .in(_U379_in),
    .clk(_U379_clk),
    .out(_U379_out)
);
assign _U380_in = _U379_out;
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign _U381_in = _U380_out;
assign _U381_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U381 (
    .in(_U381_in),
    .clk(_U381_clk),
    .out(_U381_out)
);
assign _U382_in = _U388_out;
_U382_pt__U383 _U382 (
    .in(_U382_in),
    .out(_U382_out)
);
assign _U384_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U384 (
    .in(_U384_in),
    .clk(_U384_clk),
    .out(_U384_out)
);
assign _U385_in = _U384_out;
assign _U385_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U385 (
    .in(_U385_in),
    .clk(_U385_clk),
    .out(_U385_out)
);
assign _U386_in = _U385_out;
assign _U386_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U386 (
    .in(_U386_in),
    .clk(_U386_clk),
    .out(_U386_out)
);
assign _U387_in = _U386_out;
assign _U387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U387 (
    .in(_U387_in),
    .clk(_U387_clk),
    .out(_U387_out)
);
assign _U388_in = _U387_out;
assign _U388_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U388 (
    .in(_U388_in),
    .clk(_U388_clk),
    .out(_U388_out)
);
assign _U389_in = _U395_out;
_U389_pt__U390 _U389 (
    .in(_U389_in),
    .out(_U389_out)
);
assign _U391_in = in1_hw_input_global_wrapper_stencil[6];
assign _U391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U391_in),
    .clk(_U391_clk),
    .out(_U391_out)
);
assign _U392_in = _U391_out;
assign _U392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U392_in),
    .clk(_U392_clk),
    .out(_U392_out)
);
assign _U393_in = _U392_out;
assign _U393_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U393 (
    .in(_U393_in),
    .clk(_U393_clk),
    .out(_U393_out)
);
assign _U394_in = _U393_out;
assign _U394_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U394 (
    .in(_U394_in),
    .clk(_U394_clk),
    .out(_U394_out)
);
assign _U395_in = _U394_out;
assign _U395_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U395 (
    .in(_U395_in),
    .clk(_U395_clk),
    .out(_U395_out)
);
assign _U396_in = _U403_out;
_U396_pt__U397 _U396 (
    .in(_U396_in),
    .out(_U396_out)
);
assign _U398_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = _U398_out;
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign _U400_in = _U399_out;
assign _U400_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U400 (
    .in(_U400_in),
    .clk(_U400_clk),
    .out(_U400_out)
);
assign _U401_in = _U400_out;
assign _U401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U401_in),
    .clk(_U401_clk),
    .out(_U401_out)
);
assign _U402_in = _U401_out;
assign _U402_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U402 (
    .in(_U402_in),
    .clk(_U402_clk),
    .out(_U402_out)
);
assign _U403_in = _U402_out;
assign _U403_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U403 (
    .in(_U403_in),
    .clk(_U403_clk),
    .out(_U403_out)
);
assign _U404_in = _U411_out;
_U404_pt__U405 _U404 (
    .in(_U404_in),
    .out(_U404_out)
);
assign _U406_in = in1_hw_input_global_wrapper_stencil[7];
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = _U406_out;
assign _U407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U407 (
    .in(_U407_in),
    .clk(_U407_clk),
    .out(_U407_out)
);
assign _U408_in = _U407_out;
assign _U408_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U408 (
    .in(_U408_in),
    .clk(_U408_clk),
    .out(_U408_out)
);
assign _U409_in = _U408_out;
assign _U409_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U409 (
    .in(_U409_in),
    .clk(_U409_clk),
    .out(_U409_out)
);
assign _U410_in = _U409_out;
assign _U410_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U410 (
    .in(_U410_in),
    .clk(_U410_clk),
    .out(_U410_out)
);
assign _U411_in = _U410_out;
assign _U411_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U411 (
    .in(_U411_in),
    .clk(_U411_clk),
    .out(_U411_out)
);
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U20_pt__U21 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U196_pt__U197 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U193_pt__U194 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U189_pt__U190 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U186_pt__U187 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U180_pt__U181 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U17_pt__U18 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U177_pt__U178 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U169_pt__U170 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U166_pt__U167 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U15_pt__U16 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U156_pt__U157 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U153_pt__U154 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U141_pt__U142 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U13_pt__U14 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U138_pt__U139 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U135_pt__U136 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U121_pt__U122 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U119_pt__U120 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U115_pt__U116 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U10_pt__U11 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_4_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U10_in;
wire [15:0] _U10_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U102_in;
wire _U102_clk;
wire [15:0] _U102_out;
wire [15:0] _U103_in;
wire _U103_clk;
wire [15:0] _U103_out;
wire [15:0] _U104_in;
wire _U104_clk;
wire [15:0] _U104_out;
wire [15:0] _U105_in;
wire _U105_clk;
wire [15:0] _U105_out;
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire _U108_clk;
wire [15:0] _U108_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
wire [15:0] _U110_in;
wire _U110_clk;
wire [15:0] _U110_out;
wire [15:0] _U111_in;
wire _U111_clk;
wire [15:0] _U111_out;
wire [15:0] _U112_in;
wire _U112_clk;
wire [15:0] _U112_out;
wire [15:0] _U113_in;
wire _U113_clk;
wire [15:0] _U113_out;
wire [15:0] _U114_in;
wire _U114_clk;
wire [15:0] _U114_out;
wire [15:0] _U115_in;
wire [15:0] _U115_out;
wire [15:0] _U117_in;
wire _U117_clk;
wire [15:0] _U117_out;
wire [15:0] _U118_in;
wire _U118_clk;
wire [15:0] _U118_out;
wire [15:0] _U119_in;
wire [15:0] _U12_in;
wire _U12_clk;
wire [15:0] _U12_out;
wire [15:0] _U121_in;
wire [15:0] _U121_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
wire [15:0] _U125_in;
wire _U125_clk;
wire [15:0] _U125_out;
wire [15:0] _U126_in;
wire _U126_clk;
wire [15:0] _U126_out;
wire [15:0] _U127_in;
wire _U127_clk;
wire [15:0] _U127_out;
wire [15:0] _U128_in;
wire _U128_clk;
wire [15:0] _U128_out;
wire [15:0] _U129_in;
wire _U129_clk;
wire [15:0] _U129_out;
wire [15:0] _U13_in;
wire [15:0] _U13_out;
wire [15:0] _U130_in;
wire _U130_clk;
wire [15:0] _U130_out;
wire [15:0] _U131_in;
wire _U131_clk;
wire [15:0] _U131_out;
wire [15:0] _U132_in;
wire _U132_clk;
wire [15:0] _U132_out;
wire [15:0] _U133_in;
wire _U133_clk;
wire [15:0] _U133_out;
wire [15:0] _U134_in;
wire _U134_clk;
wire [15:0] _U134_out;
wire [15:0] _U135_in;
wire [15:0] _U135_out;
wire [15:0] _U137_in;
wire _U137_clk;
wire [15:0] _U137_out;
wire [15:0] _U138_in;
wire [15:0] _U138_out;
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire [15:0] _U141_out;
wire [15:0] _U143_in;
wire _U143_clk;
wire [15:0] _U143_out;
wire [15:0] _U144_in;
wire _U144_clk;
wire [15:0] _U144_out;
wire [15:0] _U145_in;
wire _U145_clk;
wire [15:0] _U145_out;
wire [15:0] _U146_in;
wire _U146_clk;
wire [15:0] _U146_out;
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire _U148_clk;
wire [15:0] _U148_out;
wire [15:0] _U149_in;
wire _U149_clk;
wire [15:0] _U149_out;
wire [15:0] _U15_in;
wire [15:0] _U15_out;
wire [15:0] _U150_in;
wire _U150_clk;
wire [15:0] _U150_out;
wire [15:0] _U151_in;
wire _U151_clk;
wire [15:0] _U151_out;
wire [15:0] _U152_in;
wire _U152_clk;
wire [15:0] _U152_out;
wire [15:0] _U153_in;
wire [15:0] _U153_out;
wire [15:0] _U155_in;
wire _U155_clk;
wire [15:0] _U155_out;
wire [15:0] _U156_in;
wire [15:0] _U156_out;
wire [15:0] _U158_in;
wire _U158_clk;
wire [15:0] _U158_out;
wire [15:0] _U159_in;
wire _U159_clk;
wire [15:0] _U159_out;
wire [15:0] _U160_in;
wire _U160_clk;
wire [15:0] _U160_out;
wire [15:0] _U161_in;
wire _U161_clk;
wire [15:0] _U161_out;
wire [15:0] _U162_in;
wire _U162_clk;
wire [15:0] _U162_out;
wire [15:0] _U163_in;
wire _U163_clk;
wire [15:0] _U163_out;
wire [15:0] _U164_in;
wire _U164_clk;
wire [15:0] _U164_out;
wire [15:0] _U165_in;
wire _U165_clk;
wire [15:0] _U165_out;
wire [15:0] _U166_in;
wire [15:0] _U166_out;
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
wire [15:0] _U169_in;
wire [15:0] _U169_out;
wire [15:0] _U17_in;
wire [15:0] _U17_out;
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire _U172_clk;
wire [15:0] _U172_out;
wire [15:0] _U173_in;
wire _U173_clk;
wire [15:0] _U173_out;
wire [15:0] _U174_in;
wire _U174_clk;
wire [15:0] _U174_out;
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
wire [15:0] _U176_in;
wire _U176_clk;
wire [15:0] _U176_out;
wire [15:0] _U177_in;
wire [15:0] _U177_out;
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
wire [15:0] _U180_in;
wire [15:0] _U180_out;
wire [15:0] _U182_in;
wire _U182_clk;
wire [15:0] _U182_out;
wire [15:0] _U183_in;
wire _U183_clk;
wire [15:0] _U183_out;
wire [15:0] _U184_in;
wire _U184_clk;
wire [15:0] _U184_out;
wire [15:0] _U185_in;
wire _U185_clk;
wire [15:0] _U185_out;
wire [15:0] _U186_in;
wire [15:0] _U186_out;
wire [15:0] _U188_in;
wire _U188_clk;
wire [15:0] _U188_out;
wire [15:0] _U189_in;
wire [15:0] _U189_out;
wire [15:0] _U19_in;
wire _U19_clk;
wire [15:0] _U19_out;
wire [15:0] _U191_in;
wire _U191_clk;
wire [15:0] _U191_out;
wire [15:0] _U192_in;
wire _U192_clk;
wire [15:0] _U192_out;
wire [15:0] _U193_in;
wire [15:0] _U193_out;
wire [15:0] _U195_in;
wire _U195_clk;
wire [15:0] _U195_out;
wire [15:0] _U196_in;
wire [15:0] _U196_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire _U199_clk;
wire [15:0] _U199_out;
wire [15:0] _U20_in;
wire [15:0] _U20_out;
wire [15:0] _U200_in;
wire _U200_clk;
wire [15:0] _U200_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
wire [15:0] _U202_in;
wire _U202_clk;
wire [15:0] _U202_out;
wire [15:0] _U203_in;
wire _U203_clk;
wire [15:0] _U203_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U205_in;
wire _U205_clk;
wire [15:0] _U205_out;
wire [15:0] _U206_in;
wire _U206_clk;
wire [15:0] _U206_out;
wire [15:0] _U207_in;
wire _U207_clk;
wire [15:0] _U207_out;
wire [15:0] _U208_in;
wire _U208_clk;
wire [15:0] _U208_out;
wire [15:0] _U209_in;
wire _U209_clk;
wire [15:0] _U209_out;
wire [15:0] _U210_in;
wire _U210_clk;
wire [15:0] _U210_out;
wire [15:0] _U22_in;
wire _U22_clk;
wire [15:0] _U22_out;
wire [15:0] _U23_in;
wire [15:0] _U23_out;
wire [15:0] _U25_in;
wire _U25_clk;
wire [15:0] _U25_out;
wire [15:0] _U26_in;
wire _U26_clk;
wire [15:0] _U26_out;
wire [15:0] _U27_in;
wire [15:0] _U27_out;
wire [15:0] _U29_in;
wire _U29_clk;
wire [15:0] _U29_out;
wire [15:0] _U30_in;
wire _U30_clk;
wire [15:0] _U30_out;
wire [15:0] _U31_in;
wire [15:0] _U31_out;
wire [15:0] _U33_in;
wire _U33_clk;
wire [15:0] _U33_out;
wire [15:0] _U34_in;
wire _U34_clk;
wire [15:0] _U34_out;
wire [15:0] _U35_in;
wire _U35_clk;
wire [15:0] _U35_out;
wire [15:0] _U36_in;
wire [15:0] _U36_out;
wire [15:0] _U38_in;
wire _U38_clk;
wire [15:0] _U38_out;
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
wire [15:0] _U40_in;
wire _U40_clk;
wire [15:0] _U40_out;
wire [15:0] _U41_in;
wire [15:0] _U41_out;
wire [15:0] _U43_in;
wire _U43_clk;
wire [15:0] _U43_out;
wire [15:0] _U44_in;
wire _U44_clk;
wire [15:0] _U44_out;
wire [15:0] _U45_in;
wire _U45_clk;
wire [15:0] _U45_out;
wire [15:0] _U46_in;
wire _U46_clk;
wire [15:0] _U46_out;
wire [15:0] _U47_in;
wire [15:0] _U47_out;
wire [15:0] _U49_in;
wire _U49_clk;
wire [15:0] _U49_out;
wire [15:0] _U50_in;
wire _U50_clk;
wire [15:0] _U50_out;
wire [15:0] _U51_in;
wire _U51_clk;
wire [15:0] _U51_out;
wire [15:0] _U52_in;
wire _U52_clk;
wire [15:0] _U52_out;
wire [15:0] _U53_in;
wire [15:0] _U53_out;
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
wire [15:0] _U56_in;
wire _U56_clk;
wire [15:0] _U56_out;
wire [15:0] _U57_in;
wire _U57_clk;
wire [15:0] _U57_out;
wire [15:0] _U58_in;
wire _U58_clk;
wire [15:0] _U58_out;
wire [15:0] _U59_in;
wire _U59_clk;
wire [15:0] _U59_out;
wire [15:0] _U60_in;
wire [15:0] _U60_out;
wire [15:0] _U62_in;
wire _U62_clk;
wire [15:0] _U62_out;
wire [15:0] _U63_in;
wire _U63_clk;
wire [15:0] _U63_out;
wire [15:0] _U64_in;
wire _U64_clk;
wire [15:0] _U64_out;
wire [15:0] _U65_in;
wire _U65_clk;
wire [15:0] _U65_out;
wire [15:0] _U66_in;
wire _U66_clk;
wire [15:0] _U66_out;
wire [15:0] _U67_in;
wire [15:0] _U67_out;
wire [15:0] _U69_in;
wire _U69_clk;
wire [15:0] _U69_out;
wire [15:0] _U70_in;
wire _U70_clk;
wire [15:0] _U70_out;
wire [15:0] _U71_in;
wire _U71_clk;
wire [15:0] _U71_out;
wire [15:0] _U72_in;
wire _U72_clk;
wire [15:0] _U72_out;
wire [15:0] _U73_in;
wire _U73_clk;
wire [15:0] _U73_out;
wire [15:0] _U74_in;
wire _U74_clk;
wire [15:0] _U74_out;
wire [15:0] _U75_in;
wire [15:0] _U75_out;
wire [15:0] _U77_in;
wire _U77_clk;
wire [15:0] _U77_out;
wire [15:0] _U78_in;
wire _U78_clk;
wire [15:0] _U78_out;
wire [15:0] _U79_in;
wire _U79_clk;
wire [15:0] _U79_out;
wire [15:0] _U80_in;
wire _U80_clk;
wire [15:0] _U80_out;
wire [15:0] _U81_in;
wire _U81_clk;
wire [15:0] _U81_out;
wire [15:0] _U82_in;
wire _U82_clk;
wire [15:0] _U82_out;
wire [15:0] _U83_in;
wire [15:0] _U83_out;
wire [15:0] _U85_in;
wire _U85_clk;
wire [15:0] _U85_out;
wire [15:0] _U86_in;
wire _U86_clk;
wire [15:0] _U86_out;
wire [15:0] _U87_in;
wire _U87_clk;
wire [15:0] _U87_out;
wire [15:0] _U88_in;
wire _U88_clk;
wire [15:0] _U88_out;
wire [15:0] _U89_in;
wire _U89_clk;
wire [15:0] _U89_out;
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
wire [15:0] _U93_in;
wire _U93_clk;
wire [15:0] _U93_out;
wire [15:0] _U94_in;
wire _U94_clk;
wire [15:0] _U94_out;
wire [15:0] _U95_in;
wire _U95_clk;
wire [15:0] _U95_out;
wire [15:0] _U96_in;
wire _U96_clk;
wire [15:0] _U96_out;
wire [15:0] _U97_in;
wire _U97_clk;
wire [15:0] _U97_out;
wire [15:0] _U98_in;
wire _U98_clk;
wire [15:0] _U98_out;
wire [15:0] _U99_in;
wire [15:0] _U99_out;
assign _U10_in = _U12_out;
_U10_pt__U11 _U10 (
    .in(_U10_in),
    .out(_U10_out)
);
assign _U101_in = in1_hw_input_global_wrapper_stencil[7];
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U102_in = _U101_out;
assign _U102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U102_in),
    .clk(_U102_clk),
    .out(_U102_out)
);
assign _U103_in = _U102_out;
assign _U103_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U103 (
    .in(_U103_in),
    .clk(_U103_clk),
    .out(_U103_out)
);
assign _U104_in = _U103_out;
assign _U104_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U104 (
    .in(_U104_in),
    .clk(_U104_clk),
    .out(_U104_out)
);
assign _U105_in = _U104_out;
assign _U105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U105 (
    .in(_U105_in),
    .clk(_U105_clk),
    .out(_U105_out)
);
assign _U106_in = _U105_out;
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = _U106_out;
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = _U107_out;
assign _U108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U108_in),
    .clk(_U108_clk),
    .out(_U108_out)
);
assign _U109_in = _U108_out;
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign _U110_in = _U109_out;
assign _U110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U110_in),
    .clk(_U110_clk),
    .out(_U110_out)
);
assign _U111_in = _U110_out;
assign _U111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U111 (
    .in(_U111_in),
    .clk(_U111_clk),
    .out(_U111_out)
);
assign _U112_in = _U111_out;
assign _U112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U112_in),
    .clk(_U112_clk),
    .out(_U112_out)
);
assign _U113_in = _U112_out;
assign _U113_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U113 (
    .in(_U113_in),
    .clk(_U113_clk),
    .out(_U113_out)
);
assign _U114_in = _U113_out;
assign _U114_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U114 (
    .in(_U114_in),
    .clk(_U114_clk),
    .out(_U114_out)
);
assign _U115_in = _U118_out;
_U115_pt__U116 _U115 (
    .in(_U115_in),
    .out(_U115_out)
);
assign _U117_in = 16'(_U196_out + _U138_out);
assign _U117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U117 (
    .in(_U117_in),
    .clk(_U117_clk),
    .out(_U117_out)
);
assign _U118_in = _U117_out;
assign _U118_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U118 (
    .in(_U118_in),
    .clk(_U118_clk),
    .out(_U118_out)
);
assign _U119_in = 16'(_U10_out + _U115_out);
_U119_pt__U120 _U119 (
    .in(_U119_in),
    .out(out_conv_stencil)
);
assign _U12_in = 16'(_U83_out * _U99_out);
assign _U12_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U12 (
    .in(_U12_in),
    .clk(_U12_clk),
    .out(_U12_out)
);
assign _U121_in = _U134_out;
_U121_pt__U122 _U121 (
    .in(_U121_in),
    .out(_U121_out)
);
assign _U123_in = 16'(_U13_out * _U15_out);
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = _U123_out;
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign _U125_in = _U124_out;
assign _U125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U125 (
    .in(_U125_in),
    .clk(_U125_clk),
    .out(_U125_out)
);
assign _U126_in = _U125_out;
assign _U126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(_U126_in),
    .clk(_U126_clk),
    .out(_U126_out)
);
assign _U127_in = _U126_out;
assign _U127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U127_in),
    .clk(_U127_clk),
    .out(_U127_out)
);
assign _U128_in = _U127_out;
assign _U128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U128_in),
    .clk(_U128_clk),
    .out(_U128_out)
);
assign _U129_in = _U128_out;
assign _U129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U129_in),
    .clk(_U129_clk),
    .out(_U129_out)
);
assign _U13_in = in2_hw_kernel_global_wrapper_stencil[0];
_U13_pt__U14 _U13 (
    .in(_U13_in),
    .out(_U13_out)
);
assign _U130_in = _U129_out;
assign _U130_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U130 (
    .in(_U130_in),
    .clk(_U130_clk),
    .out(_U130_out)
);
assign _U131_in = _U130_out;
assign _U131_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U131 (
    .in(_U131_in),
    .clk(_U131_clk),
    .out(_U131_out)
);
assign _U132_in = _U131_out;
assign _U132_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(_U132_in),
    .clk(_U132_clk),
    .out(_U132_out)
);
assign _U133_in = _U132_out;
assign _U133_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U133 (
    .in(_U133_in),
    .clk(_U133_clk),
    .out(_U133_out)
);
assign _U134_in = _U133_out;
assign _U134_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U134 (
    .in(_U134_in),
    .clk(_U134_clk),
    .out(_U134_out)
);
assign _U135_in = _U137_out;
_U135_pt__U136 _U135 (
    .in(_U135_in),
    .out(_U135_out)
);
assign _U137_in = 16'(_U141_out + _U153_out);
assign _U137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U137 (
    .in(_U137_in),
    .clk(_U137_clk),
    .out(_U137_out)
);
assign _U138_in = _U140_out;
_U138_pt__U139 _U138 (
    .in(_U138_in),
    .out(_U138_out)
);
assign _U140_in = 16'(_U121_out + _U135_out);
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = _U152_out;
_U141_pt__U142 _U141 (
    .in(_U141_in),
    .out(_U141_out)
);
assign _U143_in = 16'(_U17_out * _U20_out);
assign _U143_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U143 (
    .in(_U143_in),
    .clk(_U143_clk),
    .out(_U143_out)
);
assign _U144_in = _U143_out;
assign _U144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U144 (
    .in(_U144_in),
    .clk(_U144_clk),
    .out(_U144_out)
);
assign _U145_in = _U144_out;
assign _U145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U145_in),
    .clk(_U145_clk),
    .out(_U145_out)
);
assign _U146_in = _U145_out;
assign _U146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U146_in),
    .clk(_U146_clk),
    .out(_U146_out)
);
assign _U147_in = _U146_out;
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = _U147_out;
assign _U148_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U148 (
    .in(_U148_in),
    .clk(_U148_clk),
    .out(_U148_out)
);
assign _U149_in = _U148_out;
assign _U149_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U149 (
    .in(_U149_in),
    .clk(_U149_clk),
    .out(_U149_out)
);
assign _U15_in = in1_hw_input_global_wrapper_stencil[0];
_U15_pt__U16 _U15 (
    .in(_U15_in),
    .out(_U15_out)
);
assign _U150_in = _U149_out;
assign _U150_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U150 (
    .in(_U150_in),
    .clk(_U150_clk),
    .out(_U150_out)
);
assign _U151_in = _U150_out;
assign _U151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(_U151_in),
    .clk(_U151_clk),
    .out(_U151_out)
);
assign _U152_in = _U151_out;
assign _U152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U152 (
    .in(_U152_in),
    .clk(_U152_clk),
    .out(_U152_out)
);
assign _U153_in = _U155_out;
_U153_pt__U154 _U153 (
    .in(_U153_in),
    .out(_U153_out)
);
assign _U155_in = 16'(_U156_out + _U166_out);
assign _U155_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U155 (
    .in(_U155_in),
    .clk(_U155_clk),
    .out(_U155_out)
);
assign _U156_in = _U165_out;
_U156_pt__U157 _U156 (
    .in(_U156_in),
    .out(_U156_out)
);
assign _U158_in = 16'(_U23_out * _U27_out);
assign _U158_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U158 (
    .in(_U158_in),
    .clk(_U158_clk),
    .out(_U158_out)
);
assign _U159_in = _U158_out;
assign _U159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U159_in),
    .clk(_U159_clk),
    .out(_U159_out)
);
assign _U160_in = _U159_out;
assign _U160_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U160 (
    .in(_U160_in),
    .clk(_U160_clk),
    .out(_U160_out)
);
assign _U161_in = _U160_out;
assign _U161_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U161 (
    .in(_U161_in),
    .clk(_U161_clk),
    .out(_U161_out)
);
assign _U162_in = _U161_out;
assign _U162_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U162 (
    .in(_U162_in),
    .clk(_U162_clk),
    .out(_U162_out)
);
assign _U163_in = _U162_out;
assign _U163_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(_U163_in),
    .clk(_U163_clk),
    .out(_U163_out)
);
assign _U164_in = _U163_out;
assign _U164_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(_U164_in),
    .clk(_U164_clk),
    .out(_U164_out)
);
assign _U165_in = _U164_out;
assign _U165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(_U165_in),
    .clk(_U165_clk),
    .out(_U165_out)
);
assign _U166_in = _U168_out;
_U166_pt__U167 _U166 (
    .in(_U166_in),
    .out(_U166_out)
);
assign _U168_in = 16'(_U169_out + _U177_out);
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign _U169_in = _U176_out;
_U169_pt__U170 _U169 (
    .in(_U169_in),
    .out(_U169_out)
);
assign _U17_in = _U19_out;
_U17_pt__U18 _U17 (
    .in(_U17_in),
    .out(_U17_out)
);
assign _U171_in = 16'(_U31_out * _U36_out);
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = _U171_out;
assign _U172_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(_U172_in),
    .clk(_U172_clk),
    .out(_U172_out)
);
assign _U173_in = _U172_out;
assign _U173_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U173 (
    .in(_U173_in),
    .clk(_U173_clk),
    .out(_U173_out)
);
assign _U174_in = _U173_out;
assign _U174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(_U174_in),
    .clk(_U174_clk),
    .out(_U174_out)
);
assign _U175_in = _U174_out;
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign _U176_in = _U175_out;
assign _U176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U176 (
    .in(_U176_in),
    .clk(_U176_clk),
    .out(_U176_out)
);
assign _U177_in = _U179_out;
_U177_pt__U178 _U177 (
    .in(_U177_in),
    .out(_U177_out)
);
assign _U179_in = 16'(_U180_out + _U186_out);
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign _U180_in = _U185_out;
_U180_pt__U181 _U180 (
    .in(_U180_in),
    .out(_U180_out)
);
assign _U182_in = 16'(_U41_out * _U47_out);
assign _U182_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U182 (
    .in(_U182_in),
    .clk(_U182_clk),
    .out(_U182_out)
);
assign _U183_in = _U182_out;
assign _U183_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U183 (
    .in(_U183_in),
    .clk(_U183_clk),
    .out(_U183_out)
);
assign _U184_in = _U183_out;
assign _U184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U184_in),
    .clk(_U184_clk),
    .out(_U184_out)
);
assign _U185_in = _U184_out;
assign _U185_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U185 (
    .in(_U185_in),
    .clk(_U185_clk),
    .out(_U185_out)
);
assign _U186_in = _U188_out;
_U186_pt__U187 _U186 (
    .in(_U186_in),
    .out(_U186_out)
);
assign _U188_in = 16'(_U189_out + _U193_out);
assign _U188_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U188 (
    .in(_U188_in),
    .clk(_U188_clk),
    .out(_U188_out)
);
assign _U189_in = _U192_out;
_U189_pt__U190 _U189 (
    .in(_U189_in),
    .out(_U189_out)
);
assign _U19_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U19_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U19 (
    .in(_U19_in),
    .clk(_U19_clk),
    .out(_U19_out)
);
assign _U191_in = 16'(_U53_out * _U60_out);
assign _U191_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U191_in),
    .clk(_U191_clk),
    .out(_U191_out)
);
assign _U192_in = _U191_out;
assign _U192_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U192_in),
    .clk(_U192_clk),
    .out(_U192_out)
);
assign _U193_in = _U195_out;
_U193_pt__U194 _U193 (
    .in(_U193_in),
    .out(_U193_out)
);
assign _U195_in = 16'(_U67_out * _U75_out);
assign _U195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U195 (
    .in(_U195_in),
    .clk(_U195_clk),
    .out(_U195_out)
);
assign _U196_in = _U210_out;
_U196_pt__U197 _U196 (
    .in(_U196_in),
    .out(_U196_out)
);
assign _U198_in = in0_conv_stencil[0];
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = _U198_out;
assign _U199_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U199 (
    .in(_U199_in),
    .clk(_U199_clk),
    .out(_U199_out)
);
assign _U20_in = _U22_out;
_U20_pt__U21 _U20 (
    .in(_U20_in),
    .out(_U20_out)
);
assign _U200_in = _U199_out;
assign _U200_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U200 (
    .in(_U200_in),
    .clk(_U200_clk),
    .out(_U200_out)
);
assign _U201_in = _U200_out;
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign _U202_in = _U201_out;
assign _U202_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U202 (
    .in(_U202_in),
    .clk(_U202_clk),
    .out(_U202_out)
);
assign _U203_in = _U202_out;
assign _U203_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U203 (
    .in(_U203_in),
    .clk(_U203_clk),
    .out(_U203_out)
);
assign _U204_in = _U203_out;
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U205_in = _U204_out;
assign _U205_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U205 (
    .in(_U205_in),
    .clk(_U205_clk),
    .out(_U205_out)
);
assign _U206_in = _U205_out;
assign _U206_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U206 (
    .in(_U206_in),
    .clk(_U206_clk),
    .out(_U206_out)
);
assign _U207_in = _U206_out;
assign _U207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(_U207_in),
    .clk(_U207_clk),
    .out(_U207_out)
);
assign _U208_in = _U207_out;
assign _U208_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U208 (
    .in(_U208_in),
    .clk(_U208_clk),
    .out(_U208_out)
);
assign _U209_in = _U208_out;
assign _U209_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U209 (
    .in(_U209_in),
    .clk(_U209_clk),
    .out(_U209_out)
);
assign _U210_in = _U209_out;
assign _U210_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U210 (
    .in(_U210_in),
    .clk(_U210_clk),
    .out(_U210_out)
);
assign _U22_in = in1_hw_input_global_wrapper_stencil[1];
assign _U22_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U22 (
    .in(_U22_in),
    .clk(_U22_clk),
    .out(_U22_out)
);
assign _U23_in = _U26_out;
_U23_pt__U24 _U23 (
    .in(_U23_in),
    .out(_U23_out)
);
assign _U25_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U25_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U25 (
    .in(_U25_in),
    .clk(_U25_clk),
    .out(_U25_out)
);
assign _U26_in = _U25_out;
assign _U26_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U26 (
    .in(_U26_in),
    .clk(_U26_clk),
    .out(_U26_out)
);
assign _U27_in = _U30_out;
_U27_pt__U28 _U27 (
    .in(_U27_in),
    .out(_U27_out)
);
assign _U29_in = in1_hw_input_global_wrapper_stencil[2];
assign _U29_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U29 (
    .in(_U29_in),
    .clk(_U29_clk),
    .out(_U29_out)
);
assign _U30_in = _U29_out;
assign _U30_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U30 (
    .in(_U30_in),
    .clk(_U30_clk),
    .out(_U30_out)
);
assign _U31_in = _U35_out;
_U31_pt__U32 _U31 (
    .in(_U31_in),
    .out(_U31_out)
);
assign _U33_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U33_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U33 (
    .in(_U33_in),
    .clk(_U33_clk),
    .out(_U33_out)
);
assign _U34_in = _U33_out;
assign _U34_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U34 (
    .in(_U34_in),
    .clk(_U34_clk),
    .out(_U34_out)
);
assign _U35_in = _U34_out;
assign _U35_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U35 (
    .in(_U35_in),
    .clk(_U35_clk),
    .out(_U35_out)
);
assign _U36_in = _U40_out;
_U36_pt__U37 _U36 (
    .in(_U36_in),
    .out(_U36_out)
);
assign _U38_in = in1_hw_input_global_wrapper_stencil[3];
assign _U38_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U38 (
    .in(_U38_in),
    .clk(_U38_clk),
    .out(_U38_out)
);
assign _U39_in = _U38_out;
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign _U40_in = _U39_out;
assign _U40_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U40 (
    .in(_U40_in),
    .clk(_U40_clk),
    .out(_U40_out)
);
assign _U41_in = _U46_out;
_U41_pt__U42 _U41 (
    .in(_U41_in),
    .out(_U41_out)
);
assign _U43_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U43_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U43 (
    .in(_U43_in),
    .clk(_U43_clk),
    .out(_U43_out)
);
assign _U44_in = _U43_out;
assign _U44_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U44 (
    .in(_U44_in),
    .clk(_U44_clk),
    .out(_U44_out)
);
assign _U45_in = _U44_out;
assign _U45_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U45 (
    .in(_U45_in),
    .clk(_U45_clk),
    .out(_U45_out)
);
assign _U46_in = _U45_out;
assign _U46_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(_U46_in),
    .clk(_U46_clk),
    .out(_U46_out)
);
assign _U47_in = _U52_out;
_U47_pt__U48 _U47 (
    .in(_U47_in),
    .out(_U47_out)
);
assign _U49_in = in1_hw_input_global_wrapper_stencil[4];
assign _U49_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U49_in),
    .clk(_U49_clk),
    .out(_U49_out)
);
assign _U50_in = _U49_out;
assign _U50_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U50 (
    .in(_U50_in),
    .clk(_U50_clk),
    .out(_U50_out)
);
assign _U51_in = _U50_out;
assign _U51_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U51 (
    .in(_U51_in),
    .clk(_U51_clk),
    .out(_U51_out)
);
assign _U52_in = _U51_out;
assign _U52_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U52 (
    .in(_U52_in),
    .clk(_U52_clk),
    .out(_U52_out)
);
assign _U53_in = _U59_out;
_U53_pt__U54 _U53 (
    .in(_U53_in),
    .out(_U53_out)
);
assign _U55_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign _U56_in = _U55_out;
assign _U56_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U56 (
    .in(_U56_in),
    .clk(_U56_clk),
    .out(_U56_out)
);
assign _U57_in = _U56_out;
assign _U57_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U57 (
    .in(_U57_in),
    .clk(_U57_clk),
    .out(_U57_out)
);
assign _U58_in = _U57_out;
assign _U58_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U58 (
    .in(_U58_in),
    .clk(_U58_clk),
    .out(_U58_out)
);
assign _U59_in = _U58_out;
assign _U59_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U59_in),
    .clk(_U59_clk),
    .out(_U59_out)
);
assign _U60_in = _U66_out;
_U60_pt__U61 _U60 (
    .in(_U60_in),
    .out(_U60_out)
);
assign _U62_in = in1_hw_input_global_wrapper_stencil[5];
assign _U62_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U62 (
    .in(_U62_in),
    .clk(_U62_clk),
    .out(_U62_out)
);
assign _U63_in = _U62_out;
assign _U63_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U63 (
    .in(_U63_in),
    .clk(_U63_clk),
    .out(_U63_out)
);
assign _U64_in = _U63_out;
assign _U64_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U64 (
    .in(_U64_in),
    .clk(_U64_clk),
    .out(_U64_out)
);
assign _U65_in = _U64_out;
assign _U65_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U65 (
    .in(_U65_in),
    .clk(_U65_clk),
    .out(_U65_out)
);
assign _U66_in = _U65_out;
assign _U66_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(_U66_in),
    .clk(_U66_clk),
    .out(_U66_out)
);
assign _U67_in = _U74_out;
_U67_pt__U68 _U67 (
    .in(_U67_in),
    .out(_U67_out)
);
assign _U69_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U69_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U69 (
    .in(_U69_in),
    .clk(_U69_clk),
    .out(_U69_out)
);
assign _U70_in = _U69_out;
assign _U70_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U70 (
    .in(_U70_in),
    .clk(_U70_clk),
    .out(_U70_out)
);
assign _U71_in = _U70_out;
assign _U71_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U71 (
    .in(_U71_in),
    .clk(_U71_clk),
    .out(_U71_out)
);
assign _U72_in = _U71_out;
assign _U72_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U72 (
    .in(_U72_in),
    .clk(_U72_clk),
    .out(_U72_out)
);
assign _U73_in = _U72_out;
assign _U73_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U73 (
    .in(_U73_in),
    .clk(_U73_clk),
    .out(_U73_out)
);
assign _U74_in = _U73_out;
assign _U74_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U74 (
    .in(_U74_in),
    .clk(_U74_clk),
    .out(_U74_out)
);
assign _U75_in = _U82_out;
_U75_pt__U76 _U75 (
    .in(_U75_in),
    .out(_U75_out)
);
assign _U77_in = in1_hw_input_global_wrapper_stencil[6];
assign _U77_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U77 (
    .in(_U77_in),
    .clk(_U77_clk),
    .out(_U77_out)
);
assign _U78_in = _U77_out;
assign _U78_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U78 (
    .in(_U78_in),
    .clk(_U78_clk),
    .out(_U78_out)
);
assign _U79_in = _U78_out;
assign _U79_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(_U79_in),
    .clk(_U79_clk),
    .out(_U79_out)
);
assign _U80_in = _U79_out;
assign _U80_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(_U80_in),
    .clk(_U80_clk),
    .out(_U80_out)
);
assign _U81_in = _U80_out;
assign _U81_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U81 (
    .in(_U81_in),
    .clk(_U81_clk),
    .out(_U81_out)
);
assign _U82_in = _U81_out;
assign _U82_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U82 (
    .in(_U82_in),
    .clk(_U82_clk),
    .out(_U82_out)
);
assign _U83_in = _U98_out;
_U83_pt__U84 _U83 (
    .in(_U83_in),
    .out(_U83_out)
);
assign _U85_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U85_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U85 (
    .in(_U85_in),
    .clk(_U85_clk),
    .out(_U85_out)
);
assign _U86_in = _U85_out;
assign _U86_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U86 (
    .in(_U86_in),
    .clk(_U86_clk),
    .out(_U86_out)
);
assign _U87_in = _U86_out;
assign _U87_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U87 (
    .in(_U87_in),
    .clk(_U87_clk),
    .out(_U87_out)
);
assign _U88_in = _U87_out;
assign _U88_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U88 (
    .in(_U88_in),
    .clk(_U88_clk),
    .out(_U88_out)
);
assign _U89_in = _U88_out;
assign _U89_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U89 (
    .in(_U89_in),
    .clk(_U89_clk),
    .out(_U89_out)
);
assign _U90_in = _U89_out;
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = _U90_out;
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = _U91_out;
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign _U93_in = _U92_out;
assign _U93_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U93_in),
    .clk(_U93_clk),
    .out(_U93_out)
);
assign _U94_in = _U93_out;
assign _U94_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U94_in),
    .clk(_U94_clk),
    .out(_U94_out)
);
assign _U95_in = _U94_out;
assign _U95_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U95 (
    .in(_U95_in),
    .clk(_U95_clk),
    .out(_U95_out)
);
assign _U96_in = _U95_out;
assign _U96_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U96 (
    .in(_U96_in),
    .clk(_U96_clk),
    .out(_U96_out)
);
assign _U97_in = _U96_out;
assign _U97_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U97 (
    .in(_U97_in),
    .clk(_U97_clk),
    .out(_U97_out)
);
assign _U98_in = _U97_out;
assign _U98_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U98 (
    .in(_U98_in),
    .clk(_U98_clk),
    .out(_U98_out)
);
assign _U99_in = _U114_out;
_U99_pt__U100 _U99 (
    .in(_U99_in),
    .out(_U99_out)
);
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U0_pt__U1 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U0_in;
assign _U0_in = in0_hw_input_stencil[0];
_U0_pt__U1 _U0 (
    .in(_U0_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U103_clk;
wire [15:0] arr__U103_in [4:0];
wire [15:0] arr__U103_out [4:0];
wire arr__U110_clk;
wire [15:0] arr__U110_in [4:0];
wire [15:0] arr__U110_out [4:0];
wire arr__U117_clk;
wire [15:0] arr__U117_in [4:0];
wire [15:0] arr__U117_out [4:0];
wire arr__U124_clk;
wire [15:0] arr__U124_in [4:0];
wire [15:0] arr__U124_out [4:0];
wire arr__U131_clk;
wire [15:0] arr__U131_in [4:0];
wire [15:0] arr__U131_out [4:0];
wire arr__U138_clk;
wire [15:0] arr__U138_in [4:0];
wire [15:0] arr__U138_out [4:0];
wire arr__U145_clk;
wire [15:0] arr__U145_in [4:0];
wire [15:0] arr__U145_out [4:0];
wire arr__U152_clk;
wire [15:0] arr__U152_in [4:0];
wire [15:0] arr__U152_out [4:0];
wire arr__U159_clk;
wire [15:0] arr__U159_in [4:0];
wire [15:0] arr__U159_out [4:0];
wire arr__U166_clk;
wire [15:0] arr__U166_in [4:0];
wire [15:0] arr__U166_out [4:0];
wire arr__U173_clk;
wire [15:0] arr__U173_in [4:0];
wire [15:0] arr__U173_out [4:0];
wire arr__U180_clk;
wire [15:0] arr__U180_in [4:0];
wire [15:0] arr__U180_out [4:0];
wire arr__U187_clk;
wire [15:0] arr__U187_in [4:0];
wire [15:0] arr__U187_out [4:0];
wire arr__U194_clk;
wire [15:0] arr__U194_in [4:0];
wire [15:0] arr__U194_out [4:0];
wire arr__U201_clk;
wire [15:0] arr__U201_in [4:0];
wire [15:0] arr__U201_out [4:0];
wire arr__U208_clk;
wire [15:0] arr__U208_in [4:0];
wire [15:0] arr__U208_out [4:0];
wire arr__U215_clk;
wire [15:0] arr__U215_in [4:0];
wire [15:0] arr__U215_out [4:0];
wire arr__U229_clk;
wire [15:0] arr__U229_in [4:0];
wire [15:0] arr__U229_out [4:0];
wire arr__U236_clk;
wire [15:0] arr__U236_in [4:0];
wire [15:0] arr__U236_out [4:0];
wire arr__U262_clk;
wire [15:0] arr__U262_in [4:0];
wire [15:0] arr__U262_out [4:0];
wire arr__U269_clk;
wire [15:0] arr__U269_in [4:0];
wire [15:0] arr__U269_out [4:0];
wire arr__U276_clk;
wire [15:0] arr__U276_in [4:0];
wire [15:0] arr__U276_out [4:0];
wire arr__U28_clk;
wire [15:0] arr__U28_in [3:0];
wire [15:0] arr__U28_out [3:0];
wire arr__U283_clk;
wire [15:0] arr__U283_in [4:0];
wire [15:0] arr__U283_out [4:0];
wire arr__U290_clk;
wire [15:0] arr__U290_in [4:0];
wire [15:0] arr__U290_out [4:0];
wire arr__U297_clk;
wire [15:0] arr__U297_in [4:0];
wire [15:0] arr__U297_out [4:0];
wire arr__U304_clk;
wire [15:0] arr__U304_in [4:0];
wire [15:0] arr__U304_out [4:0];
wire arr__U311_clk;
wire [15:0] arr__U311_in [4:0];
wire [15:0] arr__U311_out [4:0];
wire arr__U318_clk;
wire [15:0] arr__U318_in [4:0];
wire [15:0] arr__U318_out [4:0];
wire arr__U325_clk;
wire [15:0] arr__U325_in [4:0];
wire [15:0] arr__U325_out [4:0];
wire arr__U332_clk;
wire [15:0] arr__U332_in [4:0];
wire [15:0] arr__U332_out [4:0];
wire arr__U339_clk;
wire [15:0] arr__U339_in [4:0];
wire [15:0] arr__U339_out [4:0];
wire arr__U34_clk;
wire [15:0] arr__U34_in [3:0];
wire [15:0] arr__U34_out [3:0];
wire arr__U346_clk;
wire [15:0] arr__U346_in [4:0];
wire [15:0] arr__U346_out [4:0];
wire arr__U353_clk;
wire [15:0] arr__U353_in [4:0];
wire [15:0] arr__U353_out [4:0];
wire arr__U360_clk;
wire [15:0] arr__U360_in [4:0];
wire [15:0] arr__U360_out [4:0];
wire arr__U367_clk;
wire [15:0] arr__U367_in [4:0];
wire [15:0] arr__U367_out [4:0];
wire arr__U374_clk;
wire [15:0] arr__U374_in [4:0];
wire [15:0] arr__U374_out [4:0];
wire arr__U395_clk;
wire [15:0] arr__U395_in [4:0];
wire [15:0] arr__U395_out [4:0];
wire arr__U402_clk;
wire [15:0] arr__U402_in [4:0];
wire [15:0] arr__U402_out [4:0];
wire arr__U428_clk;
wire [15:0] arr__U428_in [4:0];
wire [15:0] arr__U428_out [4:0];
wire arr__U435_clk;
wire [15:0] arr__U435_in [4:0];
wire [15:0] arr__U435_out [4:0];
wire arr__U44_clk;
wire [15:0] arr__U44_in [3:0];
wire [15:0] arr__U44_out [3:0];
wire arr__U442_clk;
wire [15:0] arr__U442_in [4:0];
wire [15:0] arr__U442_out [4:0];
wire arr__U449_clk;
wire [15:0] arr__U449_in [4:0];
wire [15:0] arr__U449_out [4:0];
wire arr__U456_clk;
wire [15:0] arr__U456_in [4:0];
wire [15:0] arr__U456_out [4:0];
wire arr__U463_clk;
wire [15:0] arr__U463_in [4:0];
wire [15:0] arr__U463_out [4:0];
wire arr__U470_clk;
wire [15:0] arr__U470_in [4:0];
wire [15:0] arr__U470_out [4:0];
wire arr__U477_clk;
wire [15:0] arr__U477_in [4:0];
wire [15:0] arr__U477_out [4:0];
wire arr__U484_clk;
wire [15:0] arr__U484_in [4:0];
wire [15:0] arr__U484_out [4:0];
wire arr__U491_clk;
wire [15:0] arr__U491_in [4:0];
wire [15:0] arr__U491_out [4:0];
wire arr__U498_clk;
wire [15:0] arr__U498_in [4:0];
wire [15:0] arr__U498_out [4:0];
wire arr__U50_clk;
wire [15:0] arr__U50_in [3:0];
wire [15:0] arr__U50_out [3:0];
wire arr__U505_clk;
wire [15:0] arr__U505_in [4:0];
wire [15:0] arr__U505_out [4:0];
wire arr__U512_clk;
wire [15:0] arr__U512_in [4:0];
wire [15:0] arr__U512_out [4:0];
wire arr__U519_clk;
wire [15:0] arr__U519_in [4:0];
wire [15:0] arr__U519_out [4:0];
wire arr__U526_clk;
wire [15:0] arr__U526_in [4:0];
wire [15:0] arr__U526_out [4:0];
wire arr__U533_clk;
wire [15:0] arr__U533_in [4:0];
wire [15:0] arr__U533_out [4:0];
wire arr__U540_clk;
wire [15:0] arr__U540_in [4:0];
wire [15:0] arr__U540_out [4:0];
wire arr__U70_clk;
wire [15:0] arr__U70_in [4:0];
wire [15:0] arr__U70_out [4:0];
wire arr__U77_clk;
wire [15:0] arr__U77_in [4:0];
wire [15:0] arr__U77_out [4:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U100_clk;
wire delay_reg__U100_in;
wire delay_reg__U100_out;
wire delay_reg__U101_clk;
wire delay_reg__U101_in;
wire delay_reg__U101_out;
wire delay_reg__U226_clk;
wire delay_reg__U226_in;
wire delay_reg__U226_out;
wire delay_reg__U227_clk;
wire delay_reg__U227_in;
wire delay_reg__U227_out;
wire delay_reg__U244_clk;
wire delay_reg__U244_in;
wire delay_reg__U244_out;
wire delay_reg__U245_clk;
wire delay_reg__U245_in;
wire delay_reg__U245_out;
wire delay_reg__U246_clk;
wire delay_reg__U246_in;
wire delay_reg__U246_out;
wire delay_reg__U247_clk;
wire delay_reg__U247_in;
wire delay_reg__U247_out;
wire delay_reg__U248_clk;
wire delay_reg__U248_in;
wire delay_reg__U248_out;
wire delay_reg__U249_clk;
wire delay_reg__U249_in;
wire delay_reg__U249_out;
wire delay_reg__U25_clk;
wire delay_reg__U25_in;
wire delay_reg__U25_out;
wire delay_reg__U250_clk;
wire delay_reg__U250_in;
wire delay_reg__U250_out;
wire delay_reg__U251_clk;
wire delay_reg__U251_in;
wire delay_reg__U251_out;
wire delay_reg__U252_clk;
wire delay_reg__U252_in;
wire delay_reg__U252_out;
wire delay_reg__U253_clk;
wire delay_reg__U253_in;
wire delay_reg__U253_out;
wire delay_reg__U254_clk;
wire delay_reg__U254_in;
wire delay_reg__U254_out;
wire delay_reg__U255_clk;
wire delay_reg__U255_in;
wire delay_reg__U255_out;
wire delay_reg__U256_clk;
wire delay_reg__U256_in;
wire delay_reg__U256_out;
wire delay_reg__U257_clk;
wire delay_reg__U257_in;
wire delay_reg__U257_out;
wire delay_reg__U258_clk;
wire delay_reg__U258_in;
wire delay_reg__U258_out;
wire delay_reg__U259_clk;
wire delay_reg__U259_in;
wire delay_reg__U259_out;
wire delay_reg__U26_clk;
wire delay_reg__U26_in;
wire delay_reg__U26_out;
wire delay_reg__U260_clk;
wire delay_reg__U260_in;
wire delay_reg__U260_out;
wire delay_reg__U392_clk;
wire delay_reg__U392_in;
wire delay_reg__U392_out;
wire delay_reg__U393_clk;
wire delay_reg__U393_in;
wire delay_reg__U393_out;
wire delay_reg__U41_clk;
wire delay_reg__U41_in;
wire delay_reg__U41_out;
wire delay_reg__U410_clk;
wire delay_reg__U410_in;
wire delay_reg__U410_out;
wire delay_reg__U411_clk;
wire delay_reg__U411_in;
wire delay_reg__U411_out;
wire delay_reg__U412_clk;
wire delay_reg__U412_in;
wire delay_reg__U412_out;
wire delay_reg__U413_clk;
wire delay_reg__U413_in;
wire delay_reg__U413_out;
wire delay_reg__U414_clk;
wire delay_reg__U414_in;
wire delay_reg__U414_out;
wire delay_reg__U415_clk;
wire delay_reg__U415_in;
wire delay_reg__U415_out;
wire delay_reg__U416_clk;
wire delay_reg__U416_in;
wire delay_reg__U416_out;
wire delay_reg__U417_clk;
wire delay_reg__U417_in;
wire delay_reg__U417_out;
wire delay_reg__U418_clk;
wire delay_reg__U418_in;
wire delay_reg__U418_out;
wire delay_reg__U419_clk;
wire delay_reg__U419_in;
wire delay_reg__U419_out;
wire delay_reg__U42_clk;
wire delay_reg__U42_in;
wire delay_reg__U42_out;
wire delay_reg__U420_clk;
wire delay_reg__U420_in;
wire delay_reg__U420_out;
wire delay_reg__U421_clk;
wire delay_reg__U421_in;
wire delay_reg__U421_out;
wire delay_reg__U422_clk;
wire delay_reg__U422_in;
wire delay_reg__U422_out;
wire delay_reg__U423_clk;
wire delay_reg__U423_in;
wire delay_reg__U423_out;
wire delay_reg__U424_clk;
wire delay_reg__U424_in;
wire delay_reg__U424_out;
wire delay_reg__U425_clk;
wire delay_reg__U425_in;
wire delay_reg__U425_out;
wire delay_reg__U426_clk;
wire delay_reg__U426_in;
wire delay_reg__U426_out;
wire delay_reg__U67_clk;
wire delay_reg__U67_in;
wire delay_reg__U67_out;
wire delay_reg__U68_clk;
wire delay_reg__U68_in;
wire delay_reg__U68_out;
wire delay_reg__U85_clk;
wire delay_reg__U85_in;
wire delay_reg__U85_out;
wire delay_reg__U86_clk;
wire delay_reg__U86_in;
wire delay_reg__U86_out;
wire delay_reg__U87_clk;
wire delay_reg__U87_in;
wire delay_reg__U87_out;
wire delay_reg__U88_clk;
wire delay_reg__U88_in;
wire delay_reg__U88_out;
wire delay_reg__U89_clk;
wire delay_reg__U89_in;
wire delay_reg__U89_out;
wire delay_reg__U90_clk;
wire delay_reg__U90_in;
wire delay_reg__U90_out;
wire delay_reg__U91_clk;
wire delay_reg__U91_in;
wire delay_reg__U91_out;
wire delay_reg__U92_clk;
wire delay_reg__U92_in;
wire delay_reg__U92_out;
wire delay_reg__U93_clk;
wire delay_reg__U93_in;
wire delay_reg__U93_out;
wire delay_reg__U94_clk;
wire delay_reg__U94_in;
wire delay_reg__U94_out;
wire delay_reg__U95_clk;
wire delay_reg__U95_in;
wire delay_reg__U95_out;
wire delay_reg__U96_clk;
wire delay_reg__U96_in;
wire delay_reg__U96_out;
wire delay_reg__U97_clk;
wire delay_reg__U97_in;
wire delay_reg__U97_out;
wire delay_reg__U98_clk;
wire delay_reg__U98_in;
wire delay_reg__U98_out;
wire delay_reg__U99_clk;
wire delay_reg__U99_in;
wire delay_reg__U99_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_rst_n;
wire op_hcompute_conv_stencil_1_port_controller_flush;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_rst_n;
wire op_hcompute_conv_stencil_2_port_controller_flush;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_rst_n;
wire op_hcompute_conv_stencil_3_port_controller_flush;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_rst_n;
wire op_hcompute_conv_stencil_4_port_controller_flush;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_rst_n;
wire op_hcompute_conv_stencil_5_port_controller_flush;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_rst_n;
wire op_hcompute_conv_stencil_port_controller_flush;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_rst_n;
wire op_hcompute_hw_output_stencil_port_controller_flush;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U103_clk = clk;
assign arr__U103_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U103_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U103_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U103_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U103_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U104 arr__U103 (
    .clk(arr__U103_clk),
    .in(arr__U103_in),
    .out(arr__U103_out)
);
assign arr__U110_clk = clk;
assign arr__U110_in[4] = arr__U103_out[4];
assign arr__U110_in[3] = arr__U103_out[3];
assign arr__U110_in[2] = arr__U103_out[2];
assign arr__U110_in[1] = arr__U103_out[1];
assign arr__U110_in[0] = arr__U103_out[0];
array_delay_U111 arr__U110 (
    .clk(arr__U110_clk),
    .in(arr__U110_in),
    .out(arr__U110_out)
);
assign arr__U117_clk = clk;
assign arr__U117_in[4] = arr__U110_out[4];
assign arr__U117_in[3] = arr__U110_out[3];
assign arr__U117_in[2] = arr__U110_out[2];
assign arr__U117_in[1] = arr__U110_out[1];
assign arr__U117_in[0] = arr__U110_out[0];
array_delay_U118 arr__U117 (
    .clk(arr__U117_clk),
    .in(arr__U117_in),
    .out(arr__U117_out)
);
assign arr__U124_clk = clk;
assign arr__U124_in[4] = arr__U117_out[4];
assign arr__U124_in[3] = arr__U117_out[3];
assign arr__U124_in[2] = arr__U117_out[2];
assign arr__U124_in[1] = arr__U117_out[1];
assign arr__U124_in[0] = arr__U117_out[0];
array_delay_U125 arr__U124 (
    .clk(arr__U124_clk),
    .in(arr__U124_in),
    .out(arr__U124_out)
);
assign arr__U131_clk = clk;
assign arr__U131_in[4] = arr__U124_out[4];
assign arr__U131_in[3] = arr__U124_out[3];
assign arr__U131_in[2] = arr__U124_out[2];
assign arr__U131_in[1] = arr__U124_out[1];
assign arr__U131_in[0] = arr__U124_out[0];
array_delay_U132 arr__U131 (
    .clk(arr__U131_clk),
    .in(arr__U131_in),
    .out(arr__U131_out)
);
assign arr__U138_clk = clk;
assign arr__U138_in[4] = arr__U131_out[4];
assign arr__U138_in[3] = arr__U131_out[3];
assign arr__U138_in[2] = arr__U131_out[2];
assign arr__U138_in[1] = arr__U131_out[1];
assign arr__U138_in[0] = arr__U131_out[0];
array_delay_U139 arr__U138 (
    .clk(arr__U138_clk),
    .in(arr__U138_in),
    .out(arr__U138_out)
);
assign arr__U145_clk = clk;
assign arr__U145_in[4] = arr__U138_out[4];
assign arr__U145_in[3] = arr__U138_out[3];
assign arr__U145_in[2] = arr__U138_out[2];
assign arr__U145_in[1] = arr__U138_out[1];
assign arr__U145_in[0] = arr__U138_out[0];
array_delay_U146 arr__U145 (
    .clk(arr__U145_clk),
    .in(arr__U145_in),
    .out(arr__U145_out)
);
assign arr__U152_clk = clk;
assign arr__U152_in[4] = arr__U145_out[4];
assign arr__U152_in[3] = arr__U145_out[3];
assign arr__U152_in[2] = arr__U145_out[2];
assign arr__U152_in[1] = arr__U145_out[1];
assign arr__U152_in[0] = arr__U145_out[0];
array_delay_U153 arr__U152 (
    .clk(arr__U152_clk),
    .in(arr__U152_in),
    .out(arr__U152_out)
);
assign arr__U159_clk = clk;
assign arr__U159_in[4] = arr__U152_out[4];
assign arr__U159_in[3] = arr__U152_out[3];
assign arr__U159_in[2] = arr__U152_out[2];
assign arr__U159_in[1] = arr__U152_out[1];
assign arr__U159_in[0] = arr__U152_out[0];
array_delay_U160 arr__U159 (
    .clk(arr__U159_clk),
    .in(arr__U159_in),
    .out(arr__U159_out)
);
assign arr__U166_clk = clk;
assign arr__U166_in[4] = arr__U159_out[4];
assign arr__U166_in[3] = arr__U159_out[3];
assign arr__U166_in[2] = arr__U159_out[2];
assign arr__U166_in[1] = arr__U159_out[1];
assign arr__U166_in[0] = arr__U159_out[0];
array_delay_U167 arr__U166 (
    .clk(arr__U166_clk),
    .in(arr__U166_in),
    .out(arr__U166_out)
);
assign arr__U173_clk = clk;
assign arr__U173_in[4] = arr__U166_out[4];
assign arr__U173_in[3] = arr__U166_out[3];
assign arr__U173_in[2] = arr__U166_out[2];
assign arr__U173_in[1] = arr__U166_out[1];
assign arr__U173_in[0] = arr__U166_out[0];
array_delay_U174 arr__U173 (
    .clk(arr__U173_clk),
    .in(arr__U173_in),
    .out(arr__U173_out)
);
assign arr__U180_clk = clk;
assign arr__U180_in[4] = arr__U173_out[4];
assign arr__U180_in[3] = arr__U173_out[3];
assign arr__U180_in[2] = arr__U173_out[2];
assign arr__U180_in[1] = arr__U173_out[1];
assign arr__U180_in[0] = arr__U173_out[0];
array_delay_U181 arr__U180 (
    .clk(arr__U180_clk),
    .in(arr__U180_in),
    .out(arr__U180_out)
);
assign arr__U187_clk = clk;
assign arr__U187_in[4] = arr__U180_out[4];
assign arr__U187_in[3] = arr__U180_out[3];
assign arr__U187_in[2] = arr__U180_out[2];
assign arr__U187_in[1] = arr__U180_out[1];
assign arr__U187_in[0] = arr__U180_out[0];
array_delay_U188 arr__U187 (
    .clk(arr__U187_clk),
    .in(arr__U187_in),
    .out(arr__U187_out)
);
assign arr__U194_clk = clk;
assign arr__U194_in[4] = arr__U187_out[4];
assign arr__U194_in[3] = arr__U187_out[3];
assign arr__U194_in[2] = arr__U187_out[2];
assign arr__U194_in[1] = arr__U187_out[1];
assign arr__U194_in[0] = arr__U187_out[0];
array_delay_U195 arr__U194 (
    .clk(arr__U194_clk),
    .in(arr__U194_in),
    .out(arr__U194_out)
);
assign arr__U201_clk = clk;
assign arr__U201_in[4] = arr__U194_out[4];
assign arr__U201_in[3] = arr__U194_out[3];
assign arr__U201_in[2] = arr__U194_out[2];
assign arr__U201_in[1] = arr__U194_out[1];
assign arr__U201_in[0] = arr__U194_out[0];
array_delay_U202 arr__U201 (
    .clk(arr__U201_clk),
    .in(arr__U201_in),
    .out(arr__U201_out)
);
assign arr__U208_clk = clk;
assign arr__U208_in[4] = arr__U201_out[4];
assign arr__U208_in[3] = arr__U201_out[3];
assign arr__U208_in[2] = arr__U201_out[2];
assign arr__U208_in[1] = arr__U201_out[1];
assign arr__U208_in[0] = arr__U201_out[0];
array_delay_U209 arr__U208 (
    .clk(arr__U208_clk),
    .in(arr__U208_in),
    .out(arr__U208_out)
);
assign arr__U215_clk = clk;
assign arr__U215_in[4] = arr__U208_out[4];
assign arr__U215_in[3] = arr__U208_out[3];
assign arr__U215_in[2] = arr__U208_out[2];
assign arr__U215_in[1] = arr__U208_out[1];
assign arr__U215_in[0] = arr__U208_out[0];
array_delay_U216 arr__U215 (
    .clk(arr__U215_clk),
    .in(arr__U215_in),
    .out(arr__U215_out)
);
assign arr__U229_clk = clk;
assign arr__U229_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U229_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U229_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U229_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U229_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U230 arr__U229 (
    .clk(arr__U229_clk),
    .in(arr__U229_in),
    .out(arr__U229_out)
);
assign arr__U236_clk = clk;
assign arr__U236_in[4] = arr__U229_out[4];
assign arr__U236_in[3] = arr__U229_out[3];
assign arr__U236_in[2] = arr__U229_out[2];
assign arr__U236_in[1] = arr__U229_out[1];
assign arr__U236_in[0] = arr__U229_out[0];
array_delay_U237 arr__U236 (
    .clk(arr__U236_clk),
    .in(arr__U236_in),
    .out(arr__U236_out)
);
assign arr__U262_clk = clk;
assign arr__U262_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U262_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U262_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U262_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U262_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U263 arr__U262 (
    .clk(arr__U262_clk),
    .in(arr__U262_in),
    .out(arr__U262_out)
);
assign arr__U269_clk = clk;
assign arr__U269_in[4] = arr__U262_out[4];
assign arr__U269_in[3] = arr__U262_out[3];
assign arr__U269_in[2] = arr__U262_out[2];
assign arr__U269_in[1] = arr__U262_out[1];
assign arr__U269_in[0] = arr__U262_out[0];
array_delay_U270 arr__U269 (
    .clk(arr__U269_clk),
    .in(arr__U269_in),
    .out(arr__U269_out)
);
assign arr__U276_clk = clk;
assign arr__U276_in[4] = arr__U269_out[4];
assign arr__U276_in[3] = arr__U269_out[3];
assign arr__U276_in[2] = arr__U269_out[2];
assign arr__U276_in[1] = arr__U269_out[1];
assign arr__U276_in[0] = arr__U269_out[0];
array_delay_U277 arr__U276 (
    .clk(arr__U276_clk),
    .in(arr__U276_in),
    .out(arr__U276_out)
);
assign arr__U28_clk = clk;
assign arr__U28_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U28_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U28_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U28_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U29 arr__U28 (
    .clk(arr__U28_clk),
    .in(arr__U28_in),
    .out(arr__U28_out)
);
assign arr__U283_clk = clk;
assign arr__U283_in[4] = arr__U276_out[4];
assign arr__U283_in[3] = arr__U276_out[3];
assign arr__U283_in[2] = arr__U276_out[2];
assign arr__U283_in[1] = arr__U276_out[1];
assign arr__U283_in[0] = arr__U276_out[0];
array_delay_U284 arr__U283 (
    .clk(arr__U283_clk),
    .in(arr__U283_in),
    .out(arr__U283_out)
);
assign arr__U290_clk = clk;
assign arr__U290_in[4] = arr__U283_out[4];
assign arr__U290_in[3] = arr__U283_out[3];
assign arr__U290_in[2] = arr__U283_out[2];
assign arr__U290_in[1] = arr__U283_out[1];
assign arr__U290_in[0] = arr__U283_out[0];
array_delay_U291 arr__U290 (
    .clk(arr__U290_clk),
    .in(arr__U290_in),
    .out(arr__U290_out)
);
assign arr__U297_clk = clk;
assign arr__U297_in[4] = arr__U290_out[4];
assign arr__U297_in[3] = arr__U290_out[3];
assign arr__U297_in[2] = arr__U290_out[2];
assign arr__U297_in[1] = arr__U290_out[1];
assign arr__U297_in[0] = arr__U290_out[0];
array_delay_U298 arr__U297 (
    .clk(arr__U297_clk),
    .in(arr__U297_in),
    .out(arr__U297_out)
);
assign arr__U304_clk = clk;
assign arr__U304_in[4] = arr__U297_out[4];
assign arr__U304_in[3] = arr__U297_out[3];
assign arr__U304_in[2] = arr__U297_out[2];
assign arr__U304_in[1] = arr__U297_out[1];
assign arr__U304_in[0] = arr__U297_out[0];
array_delay_U305 arr__U304 (
    .clk(arr__U304_clk),
    .in(arr__U304_in),
    .out(arr__U304_out)
);
assign arr__U311_clk = clk;
assign arr__U311_in[4] = arr__U304_out[4];
assign arr__U311_in[3] = arr__U304_out[3];
assign arr__U311_in[2] = arr__U304_out[2];
assign arr__U311_in[1] = arr__U304_out[1];
assign arr__U311_in[0] = arr__U304_out[0];
array_delay_U312 arr__U311 (
    .clk(arr__U311_clk),
    .in(arr__U311_in),
    .out(arr__U311_out)
);
assign arr__U318_clk = clk;
assign arr__U318_in[4] = arr__U311_out[4];
assign arr__U318_in[3] = arr__U311_out[3];
assign arr__U318_in[2] = arr__U311_out[2];
assign arr__U318_in[1] = arr__U311_out[1];
assign arr__U318_in[0] = arr__U311_out[0];
array_delay_U319 arr__U318 (
    .clk(arr__U318_clk),
    .in(arr__U318_in),
    .out(arr__U318_out)
);
assign arr__U325_clk = clk;
assign arr__U325_in[4] = arr__U318_out[4];
assign arr__U325_in[3] = arr__U318_out[3];
assign arr__U325_in[2] = arr__U318_out[2];
assign arr__U325_in[1] = arr__U318_out[1];
assign arr__U325_in[0] = arr__U318_out[0];
array_delay_U326 arr__U325 (
    .clk(arr__U325_clk),
    .in(arr__U325_in),
    .out(arr__U325_out)
);
assign arr__U332_clk = clk;
assign arr__U332_in[4] = arr__U325_out[4];
assign arr__U332_in[3] = arr__U325_out[3];
assign arr__U332_in[2] = arr__U325_out[2];
assign arr__U332_in[1] = arr__U325_out[1];
assign arr__U332_in[0] = arr__U325_out[0];
array_delay_U333 arr__U332 (
    .clk(arr__U332_clk),
    .in(arr__U332_in),
    .out(arr__U332_out)
);
assign arr__U339_clk = clk;
assign arr__U339_in[4] = arr__U332_out[4];
assign arr__U339_in[3] = arr__U332_out[3];
assign arr__U339_in[2] = arr__U332_out[2];
assign arr__U339_in[1] = arr__U332_out[1];
assign arr__U339_in[0] = arr__U332_out[0];
array_delay_U340 arr__U339 (
    .clk(arr__U339_clk),
    .in(arr__U339_in),
    .out(arr__U339_out)
);
assign arr__U34_clk = clk;
assign arr__U34_in[3] = arr__U28_out[3];
assign arr__U34_in[2] = arr__U28_out[2];
assign arr__U34_in[1] = arr__U28_out[1];
assign arr__U34_in[0] = arr__U28_out[0];
array_delay_U35 arr__U34 (
    .clk(arr__U34_clk),
    .in(arr__U34_in),
    .out(arr__U34_out)
);
assign arr__U346_clk = clk;
assign arr__U346_in[4] = arr__U339_out[4];
assign arr__U346_in[3] = arr__U339_out[3];
assign arr__U346_in[2] = arr__U339_out[2];
assign arr__U346_in[1] = arr__U339_out[1];
assign arr__U346_in[0] = arr__U339_out[0];
array_delay_U347 arr__U346 (
    .clk(arr__U346_clk),
    .in(arr__U346_in),
    .out(arr__U346_out)
);
assign arr__U353_clk = clk;
assign arr__U353_in[4] = arr__U346_out[4];
assign arr__U353_in[3] = arr__U346_out[3];
assign arr__U353_in[2] = arr__U346_out[2];
assign arr__U353_in[1] = arr__U346_out[1];
assign arr__U353_in[0] = arr__U346_out[0];
array_delay_U354 arr__U353 (
    .clk(arr__U353_clk),
    .in(arr__U353_in),
    .out(arr__U353_out)
);
assign arr__U360_clk = clk;
assign arr__U360_in[4] = arr__U353_out[4];
assign arr__U360_in[3] = arr__U353_out[3];
assign arr__U360_in[2] = arr__U353_out[2];
assign arr__U360_in[1] = arr__U353_out[1];
assign arr__U360_in[0] = arr__U353_out[0];
array_delay_U361 arr__U360 (
    .clk(arr__U360_clk),
    .in(arr__U360_in),
    .out(arr__U360_out)
);
assign arr__U367_clk = clk;
assign arr__U367_in[4] = arr__U360_out[4];
assign arr__U367_in[3] = arr__U360_out[3];
assign arr__U367_in[2] = arr__U360_out[2];
assign arr__U367_in[1] = arr__U360_out[1];
assign arr__U367_in[0] = arr__U360_out[0];
array_delay_U368 arr__U367 (
    .clk(arr__U367_clk),
    .in(arr__U367_in),
    .out(arr__U367_out)
);
assign arr__U374_clk = clk;
assign arr__U374_in[4] = arr__U367_out[4];
assign arr__U374_in[3] = arr__U367_out[3];
assign arr__U374_in[2] = arr__U367_out[2];
assign arr__U374_in[1] = arr__U367_out[1];
assign arr__U374_in[0] = arr__U367_out[0];
array_delay_U375 arr__U374 (
    .clk(arr__U374_clk),
    .in(arr__U374_in),
    .out(arr__U374_out)
);
assign arr__U395_clk = clk;
assign arr__U395_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U395_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U395_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U395_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U395_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U396 arr__U395 (
    .clk(arr__U395_clk),
    .in(arr__U395_in),
    .out(arr__U395_out)
);
assign arr__U402_clk = clk;
assign arr__U402_in[4] = arr__U395_out[4];
assign arr__U402_in[3] = arr__U395_out[3];
assign arr__U402_in[2] = arr__U395_out[2];
assign arr__U402_in[1] = arr__U395_out[1];
assign arr__U402_in[0] = arr__U395_out[0];
array_delay_U403 arr__U402 (
    .clk(arr__U402_clk),
    .in(arr__U402_in),
    .out(arr__U402_out)
);
assign arr__U428_clk = clk;
assign arr__U428_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U428_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U428_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U428_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U428_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U429 arr__U428 (
    .clk(arr__U428_clk),
    .in(arr__U428_in),
    .out(arr__U428_out)
);
assign arr__U435_clk = clk;
assign arr__U435_in[4] = arr__U428_out[4];
assign arr__U435_in[3] = arr__U428_out[3];
assign arr__U435_in[2] = arr__U428_out[2];
assign arr__U435_in[1] = arr__U428_out[1];
assign arr__U435_in[0] = arr__U428_out[0];
array_delay_U436 arr__U435 (
    .clk(arr__U435_clk),
    .in(arr__U435_in),
    .out(arr__U435_out)
);
assign arr__U44_clk = clk;
assign arr__U44_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U44_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U44_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U44_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U45 arr__U44 (
    .clk(arr__U44_clk),
    .in(arr__U44_in),
    .out(arr__U44_out)
);
assign arr__U442_clk = clk;
assign arr__U442_in[4] = arr__U435_out[4];
assign arr__U442_in[3] = arr__U435_out[3];
assign arr__U442_in[2] = arr__U435_out[2];
assign arr__U442_in[1] = arr__U435_out[1];
assign arr__U442_in[0] = arr__U435_out[0];
array_delay_U443 arr__U442 (
    .clk(arr__U442_clk),
    .in(arr__U442_in),
    .out(arr__U442_out)
);
assign arr__U449_clk = clk;
assign arr__U449_in[4] = arr__U442_out[4];
assign arr__U449_in[3] = arr__U442_out[3];
assign arr__U449_in[2] = arr__U442_out[2];
assign arr__U449_in[1] = arr__U442_out[1];
assign arr__U449_in[0] = arr__U442_out[0];
array_delay_U450 arr__U449 (
    .clk(arr__U449_clk),
    .in(arr__U449_in),
    .out(arr__U449_out)
);
assign arr__U456_clk = clk;
assign arr__U456_in[4] = arr__U449_out[4];
assign arr__U456_in[3] = arr__U449_out[3];
assign arr__U456_in[2] = arr__U449_out[2];
assign arr__U456_in[1] = arr__U449_out[1];
assign arr__U456_in[0] = arr__U449_out[0];
array_delay_U457 arr__U456 (
    .clk(arr__U456_clk),
    .in(arr__U456_in),
    .out(arr__U456_out)
);
assign arr__U463_clk = clk;
assign arr__U463_in[4] = arr__U456_out[4];
assign arr__U463_in[3] = arr__U456_out[3];
assign arr__U463_in[2] = arr__U456_out[2];
assign arr__U463_in[1] = arr__U456_out[1];
assign arr__U463_in[0] = arr__U456_out[0];
array_delay_U464 arr__U463 (
    .clk(arr__U463_clk),
    .in(arr__U463_in),
    .out(arr__U463_out)
);
assign arr__U470_clk = clk;
assign arr__U470_in[4] = arr__U463_out[4];
assign arr__U470_in[3] = arr__U463_out[3];
assign arr__U470_in[2] = arr__U463_out[2];
assign arr__U470_in[1] = arr__U463_out[1];
assign arr__U470_in[0] = arr__U463_out[0];
array_delay_U471 arr__U470 (
    .clk(arr__U470_clk),
    .in(arr__U470_in),
    .out(arr__U470_out)
);
assign arr__U477_clk = clk;
assign arr__U477_in[4] = arr__U470_out[4];
assign arr__U477_in[3] = arr__U470_out[3];
assign arr__U477_in[2] = arr__U470_out[2];
assign arr__U477_in[1] = arr__U470_out[1];
assign arr__U477_in[0] = arr__U470_out[0];
array_delay_U478 arr__U477 (
    .clk(arr__U477_clk),
    .in(arr__U477_in),
    .out(arr__U477_out)
);
assign arr__U484_clk = clk;
assign arr__U484_in[4] = arr__U477_out[4];
assign arr__U484_in[3] = arr__U477_out[3];
assign arr__U484_in[2] = arr__U477_out[2];
assign arr__U484_in[1] = arr__U477_out[1];
assign arr__U484_in[0] = arr__U477_out[0];
array_delay_U485 arr__U484 (
    .clk(arr__U484_clk),
    .in(arr__U484_in),
    .out(arr__U484_out)
);
assign arr__U491_clk = clk;
assign arr__U491_in[4] = arr__U484_out[4];
assign arr__U491_in[3] = arr__U484_out[3];
assign arr__U491_in[2] = arr__U484_out[2];
assign arr__U491_in[1] = arr__U484_out[1];
assign arr__U491_in[0] = arr__U484_out[0];
array_delay_U492 arr__U491 (
    .clk(arr__U491_clk),
    .in(arr__U491_in),
    .out(arr__U491_out)
);
assign arr__U498_clk = clk;
assign arr__U498_in[4] = arr__U491_out[4];
assign arr__U498_in[3] = arr__U491_out[3];
assign arr__U498_in[2] = arr__U491_out[2];
assign arr__U498_in[1] = arr__U491_out[1];
assign arr__U498_in[0] = arr__U491_out[0];
array_delay_U499 arr__U498 (
    .clk(arr__U498_clk),
    .in(arr__U498_in),
    .out(arr__U498_out)
);
assign arr__U50_clk = clk;
assign arr__U50_in[3] = arr__U44_out[3];
assign arr__U50_in[2] = arr__U44_out[2];
assign arr__U50_in[1] = arr__U44_out[1];
assign arr__U50_in[0] = arr__U44_out[0];
array_delay_U51 arr__U50 (
    .clk(arr__U50_clk),
    .in(arr__U50_in),
    .out(arr__U50_out)
);
assign arr__U505_clk = clk;
assign arr__U505_in[4] = arr__U498_out[4];
assign arr__U505_in[3] = arr__U498_out[3];
assign arr__U505_in[2] = arr__U498_out[2];
assign arr__U505_in[1] = arr__U498_out[1];
assign arr__U505_in[0] = arr__U498_out[0];
array_delay_U506 arr__U505 (
    .clk(arr__U505_clk),
    .in(arr__U505_in),
    .out(arr__U505_out)
);
assign arr__U512_clk = clk;
assign arr__U512_in[4] = arr__U505_out[4];
assign arr__U512_in[3] = arr__U505_out[3];
assign arr__U512_in[2] = arr__U505_out[2];
assign arr__U512_in[1] = arr__U505_out[1];
assign arr__U512_in[0] = arr__U505_out[0];
array_delay_U513 arr__U512 (
    .clk(arr__U512_clk),
    .in(arr__U512_in),
    .out(arr__U512_out)
);
assign arr__U519_clk = clk;
assign arr__U519_in[4] = arr__U512_out[4];
assign arr__U519_in[3] = arr__U512_out[3];
assign arr__U519_in[2] = arr__U512_out[2];
assign arr__U519_in[1] = arr__U512_out[1];
assign arr__U519_in[0] = arr__U512_out[0];
array_delay_U520 arr__U519 (
    .clk(arr__U519_clk),
    .in(arr__U519_in),
    .out(arr__U519_out)
);
assign arr__U526_clk = clk;
assign arr__U526_in[4] = arr__U519_out[4];
assign arr__U526_in[3] = arr__U519_out[3];
assign arr__U526_in[2] = arr__U519_out[2];
assign arr__U526_in[1] = arr__U519_out[1];
assign arr__U526_in[0] = arr__U519_out[0];
array_delay_U527 arr__U526 (
    .clk(arr__U526_clk),
    .in(arr__U526_in),
    .out(arr__U526_out)
);
assign arr__U533_clk = clk;
assign arr__U533_in[4] = arr__U526_out[4];
assign arr__U533_in[3] = arr__U526_out[3];
assign arr__U533_in[2] = arr__U526_out[2];
assign arr__U533_in[1] = arr__U526_out[1];
assign arr__U533_in[0] = arr__U526_out[0];
array_delay_U534 arr__U533 (
    .clk(arr__U533_clk),
    .in(arr__U533_in),
    .out(arr__U533_out)
);
assign arr__U540_clk = clk;
assign arr__U540_in[4] = arr__U533_out[4];
assign arr__U540_in[3] = arr__U533_out[3];
assign arr__U540_in[2] = arr__U533_out[2];
assign arr__U540_in[1] = arr__U533_out[1];
assign arr__U540_in[0] = arr__U533_out[0];
array_delay_U541 arr__U540 (
    .clk(arr__U540_clk),
    .in(arr__U540_in),
    .out(arr__U540_out)
);
assign arr__U70_clk = clk;
assign arr__U70_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U70_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U70_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U70_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U70_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U71 arr__U70 (
    .clk(arr__U70_clk),
    .in(arr__U70_in),
    .out(arr__U70_out)
);
assign arr__U77_clk = clk;
assign arr__U77_in[4] = arr__U70_out[4];
assign arr__U77_in[3] = arr__U70_out[3];
assign arr__U77_in[2] = arr__U70_out[2];
assign arr__U77_in[1] = arr__U70_out[1];
assign arr__U77_in[0] = arr__U70_out[0];
array_delay_U78 arr__U77 (
    .clk(arr__U77_clk),
    .in(arr__U77_in),
    .out(arr__U77_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U100_clk = clk;
assign delay_reg__U100_in = delay_reg__U99_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U100 (
    .clk(delay_reg__U100_clk),
    .in(delay_reg__U100_in),
    .out(delay_reg__U100_out)
);
assign delay_reg__U101_clk = clk;
assign delay_reg__U101_in = delay_reg__U100_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U101 (
    .clk(delay_reg__U101_clk),
    .in(delay_reg__U101_in),
    .out(delay_reg__U101_out)
);
assign delay_reg__U226_clk = clk;
assign delay_reg__U226_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U226 (
    .clk(delay_reg__U226_clk),
    .in(delay_reg__U226_in),
    .out(delay_reg__U226_out)
);
assign delay_reg__U227_clk = clk;
assign delay_reg__U227_in = delay_reg__U226_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U227 (
    .clk(delay_reg__U227_clk),
    .in(delay_reg__U227_in),
    .out(delay_reg__U227_out)
);
assign delay_reg__U244_clk = clk;
assign delay_reg__U244_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U244 (
    .clk(delay_reg__U244_clk),
    .in(delay_reg__U244_in),
    .out(delay_reg__U244_out)
);
assign delay_reg__U245_clk = clk;
assign delay_reg__U245_in = delay_reg__U244_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U245 (
    .clk(delay_reg__U245_clk),
    .in(delay_reg__U245_in),
    .out(delay_reg__U245_out)
);
assign delay_reg__U246_clk = clk;
assign delay_reg__U246_in = delay_reg__U245_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U246 (
    .clk(delay_reg__U246_clk),
    .in(delay_reg__U246_in),
    .out(delay_reg__U246_out)
);
assign delay_reg__U247_clk = clk;
assign delay_reg__U247_in = delay_reg__U246_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U247 (
    .clk(delay_reg__U247_clk),
    .in(delay_reg__U247_in),
    .out(delay_reg__U247_out)
);
assign delay_reg__U248_clk = clk;
assign delay_reg__U248_in = delay_reg__U247_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U248 (
    .clk(delay_reg__U248_clk),
    .in(delay_reg__U248_in),
    .out(delay_reg__U248_out)
);
assign delay_reg__U249_clk = clk;
assign delay_reg__U249_in = delay_reg__U248_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U249 (
    .clk(delay_reg__U249_clk),
    .in(delay_reg__U249_in),
    .out(delay_reg__U249_out)
);
assign delay_reg__U25_clk = clk;
assign delay_reg__U25_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U25 (
    .clk(delay_reg__U25_clk),
    .in(delay_reg__U25_in),
    .out(delay_reg__U25_out)
);
assign delay_reg__U250_clk = clk;
assign delay_reg__U250_in = delay_reg__U249_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U250 (
    .clk(delay_reg__U250_clk),
    .in(delay_reg__U250_in),
    .out(delay_reg__U250_out)
);
assign delay_reg__U251_clk = clk;
assign delay_reg__U251_in = delay_reg__U250_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U251 (
    .clk(delay_reg__U251_clk),
    .in(delay_reg__U251_in),
    .out(delay_reg__U251_out)
);
assign delay_reg__U252_clk = clk;
assign delay_reg__U252_in = delay_reg__U251_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U252 (
    .clk(delay_reg__U252_clk),
    .in(delay_reg__U252_in),
    .out(delay_reg__U252_out)
);
assign delay_reg__U253_clk = clk;
assign delay_reg__U253_in = delay_reg__U252_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U253 (
    .clk(delay_reg__U253_clk),
    .in(delay_reg__U253_in),
    .out(delay_reg__U253_out)
);
assign delay_reg__U254_clk = clk;
assign delay_reg__U254_in = delay_reg__U253_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U254 (
    .clk(delay_reg__U254_clk),
    .in(delay_reg__U254_in),
    .out(delay_reg__U254_out)
);
assign delay_reg__U255_clk = clk;
assign delay_reg__U255_in = delay_reg__U254_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U255 (
    .clk(delay_reg__U255_clk),
    .in(delay_reg__U255_in),
    .out(delay_reg__U255_out)
);
assign delay_reg__U256_clk = clk;
assign delay_reg__U256_in = delay_reg__U255_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U256 (
    .clk(delay_reg__U256_clk),
    .in(delay_reg__U256_in),
    .out(delay_reg__U256_out)
);
assign delay_reg__U257_clk = clk;
assign delay_reg__U257_in = delay_reg__U256_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U257 (
    .clk(delay_reg__U257_clk),
    .in(delay_reg__U257_in),
    .out(delay_reg__U257_out)
);
assign delay_reg__U258_clk = clk;
assign delay_reg__U258_in = delay_reg__U257_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U258 (
    .clk(delay_reg__U258_clk),
    .in(delay_reg__U258_in),
    .out(delay_reg__U258_out)
);
assign delay_reg__U259_clk = clk;
assign delay_reg__U259_in = delay_reg__U258_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U259 (
    .clk(delay_reg__U259_clk),
    .in(delay_reg__U259_in),
    .out(delay_reg__U259_out)
);
assign delay_reg__U26_clk = clk;
assign delay_reg__U26_in = delay_reg__U25_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U26 (
    .clk(delay_reg__U26_clk),
    .in(delay_reg__U26_in),
    .out(delay_reg__U26_out)
);
assign delay_reg__U260_clk = clk;
assign delay_reg__U260_in = delay_reg__U259_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U260 (
    .clk(delay_reg__U260_clk),
    .in(delay_reg__U260_in),
    .out(delay_reg__U260_out)
);
assign delay_reg__U392_clk = clk;
assign delay_reg__U392_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U392 (
    .clk(delay_reg__U392_clk),
    .in(delay_reg__U392_in),
    .out(delay_reg__U392_out)
);
assign delay_reg__U393_clk = clk;
assign delay_reg__U393_in = delay_reg__U392_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U393 (
    .clk(delay_reg__U393_clk),
    .in(delay_reg__U393_in),
    .out(delay_reg__U393_out)
);
assign delay_reg__U41_clk = clk;
assign delay_reg__U41_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U41 (
    .clk(delay_reg__U41_clk),
    .in(delay_reg__U41_in),
    .out(delay_reg__U41_out)
);
assign delay_reg__U410_clk = clk;
assign delay_reg__U410_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U410 (
    .clk(delay_reg__U410_clk),
    .in(delay_reg__U410_in),
    .out(delay_reg__U410_out)
);
assign delay_reg__U411_clk = clk;
assign delay_reg__U411_in = delay_reg__U410_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U411 (
    .clk(delay_reg__U411_clk),
    .in(delay_reg__U411_in),
    .out(delay_reg__U411_out)
);
assign delay_reg__U412_clk = clk;
assign delay_reg__U412_in = delay_reg__U411_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U412 (
    .clk(delay_reg__U412_clk),
    .in(delay_reg__U412_in),
    .out(delay_reg__U412_out)
);
assign delay_reg__U413_clk = clk;
assign delay_reg__U413_in = delay_reg__U412_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U413 (
    .clk(delay_reg__U413_clk),
    .in(delay_reg__U413_in),
    .out(delay_reg__U413_out)
);
assign delay_reg__U414_clk = clk;
assign delay_reg__U414_in = delay_reg__U413_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U414 (
    .clk(delay_reg__U414_clk),
    .in(delay_reg__U414_in),
    .out(delay_reg__U414_out)
);
assign delay_reg__U415_clk = clk;
assign delay_reg__U415_in = delay_reg__U414_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U415 (
    .clk(delay_reg__U415_clk),
    .in(delay_reg__U415_in),
    .out(delay_reg__U415_out)
);
assign delay_reg__U416_clk = clk;
assign delay_reg__U416_in = delay_reg__U415_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U416 (
    .clk(delay_reg__U416_clk),
    .in(delay_reg__U416_in),
    .out(delay_reg__U416_out)
);
assign delay_reg__U417_clk = clk;
assign delay_reg__U417_in = delay_reg__U416_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U417 (
    .clk(delay_reg__U417_clk),
    .in(delay_reg__U417_in),
    .out(delay_reg__U417_out)
);
assign delay_reg__U418_clk = clk;
assign delay_reg__U418_in = delay_reg__U417_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U418 (
    .clk(delay_reg__U418_clk),
    .in(delay_reg__U418_in),
    .out(delay_reg__U418_out)
);
assign delay_reg__U419_clk = clk;
assign delay_reg__U419_in = delay_reg__U418_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U419 (
    .clk(delay_reg__U419_clk),
    .in(delay_reg__U419_in),
    .out(delay_reg__U419_out)
);
assign delay_reg__U42_clk = clk;
assign delay_reg__U42_in = delay_reg__U41_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U42 (
    .clk(delay_reg__U42_clk),
    .in(delay_reg__U42_in),
    .out(delay_reg__U42_out)
);
assign delay_reg__U420_clk = clk;
assign delay_reg__U420_in = delay_reg__U419_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U420 (
    .clk(delay_reg__U420_clk),
    .in(delay_reg__U420_in),
    .out(delay_reg__U420_out)
);
assign delay_reg__U421_clk = clk;
assign delay_reg__U421_in = delay_reg__U420_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U421 (
    .clk(delay_reg__U421_clk),
    .in(delay_reg__U421_in),
    .out(delay_reg__U421_out)
);
assign delay_reg__U422_clk = clk;
assign delay_reg__U422_in = delay_reg__U421_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U422 (
    .clk(delay_reg__U422_clk),
    .in(delay_reg__U422_in),
    .out(delay_reg__U422_out)
);
assign delay_reg__U423_clk = clk;
assign delay_reg__U423_in = delay_reg__U422_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U423 (
    .clk(delay_reg__U423_clk),
    .in(delay_reg__U423_in),
    .out(delay_reg__U423_out)
);
assign delay_reg__U424_clk = clk;
assign delay_reg__U424_in = delay_reg__U423_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U424 (
    .clk(delay_reg__U424_clk),
    .in(delay_reg__U424_in),
    .out(delay_reg__U424_out)
);
assign delay_reg__U425_clk = clk;
assign delay_reg__U425_in = delay_reg__U424_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U425 (
    .clk(delay_reg__U425_clk),
    .in(delay_reg__U425_in),
    .out(delay_reg__U425_out)
);
assign delay_reg__U426_clk = clk;
assign delay_reg__U426_in = delay_reg__U425_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U426 (
    .clk(delay_reg__U426_clk),
    .in(delay_reg__U426_in),
    .out(delay_reg__U426_out)
);
assign delay_reg__U67_clk = clk;
assign delay_reg__U67_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U67 (
    .clk(delay_reg__U67_clk),
    .in(delay_reg__U67_in),
    .out(delay_reg__U67_out)
);
assign delay_reg__U68_clk = clk;
assign delay_reg__U68_in = delay_reg__U67_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U68 (
    .clk(delay_reg__U68_clk),
    .in(delay_reg__U68_in),
    .out(delay_reg__U68_out)
);
assign delay_reg__U85_clk = clk;
assign delay_reg__U85_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U85 (
    .clk(delay_reg__U85_clk),
    .in(delay_reg__U85_in),
    .out(delay_reg__U85_out)
);
assign delay_reg__U86_clk = clk;
assign delay_reg__U86_in = delay_reg__U85_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U86 (
    .clk(delay_reg__U86_clk),
    .in(delay_reg__U86_in),
    .out(delay_reg__U86_out)
);
assign delay_reg__U87_clk = clk;
assign delay_reg__U87_in = delay_reg__U86_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U87 (
    .clk(delay_reg__U87_clk),
    .in(delay_reg__U87_in),
    .out(delay_reg__U87_out)
);
assign delay_reg__U88_clk = clk;
assign delay_reg__U88_in = delay_reg__U87_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U88 (
    .clk(delay_reg__U88_clk),
    .in(delay_reg__U88_in),
    .out(delay_reg__U88_out)
);
assign delay_reg__U89_clk = clk;
assign delay_reg__U89_in = delay_reg__U88_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U89 (
    .clk(delay_reg__U89_clk),
    .in(delay_reg__U89_in),
    .out(delay_reg__U89_out)
);
assign delay_reg__U90_clk = clk;
assign delay_reg__U90_in = delay_reg__U89_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U90 (
    .clk(delay_reg__U90_clk),
    .in(delay_reg__U90_in),
    .out(delay_reg__U90_out)
);
assign delay_reg__U91_clk = clk;
assign delay_reg__U91_in = delay_reg__U90_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U91 (
    .clk(delay_reg__U91_clk),
    .in(delay_reg__U91_in),
    .out(delay_reg__U91_out)
);
assign delay_reg__U92_clk = clk;
assign delay_reg__U92_in = delay_reg__U91_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U92 (
    .clk(delay_reg__U92_clk),
    .in(delay_reg__U92_in),
    .out(delay_reg__U92_out)
);
assign delay_reg__U93_clk = clk;
assign delay_reg__U93_in = delay_reg__U92_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U93 (
    .clk(delay_reg__U93_clk),
    .in(delay_reg__U93_in),
    .out(delay_reg__U93_out)
);
assign delay_reg__U94_clk = clk;
assign delay_reg__U94_in = delay_reg__U93_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U94 (
    .clk(delay_reg__U94_clk),
    .in(delay_reg__U94_in),
    .out(delay_reg__U94_out)
);
assign delay_reg__U95_clk = clk;
assign delay_reg__U95_in = delay_reg__U94_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U95 (
    .clk(delay_reg__U95_clk),
    .in(delay_reg__U95_in),
    .out(delay_reg__U95_out)
);
assign delay_reg__U96_clk = clk;
assign delay_reg__U96_in = delay_reg__U95_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U96 (
    .clk(delay_reg__U96_clk),
    .in(delay_reg__U96_in),
    .out(delay_reg__U96_out)
);
assign delay_reg__U97_clk = clk;
assign delay_reg__U97_in = delay_reg__U96_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U97 (
    .clk(delay_reg__U97_clk),
    .in(delay_reg__U97_in),
    .out(delay_reg__U97_out)
);
assign delay_reg__U98_clk = clk;
assign delay_reg__U98_in = delay_reg__U97_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U98 (
    .clk(delay_reg__U98_clk),
    .in(delay_reg__U98_in),
    .out(delay_reg__U98_out)
);
assign delay_reg__U99_clk = clk;
assign delay_reg__U99_in = delay_reg__U98_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U99 (
    .clk(delay_reg__U99_clk),
    .in(delay_reg__U99_in),
    .out(delay_reg__U99_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U10 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U11 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
assign op_hcompute_conv_stencil_1_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_1_port_controller_flush = flush;
affine_controller__U7 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_1_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_1_port_controller_flush),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U8 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U9 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U12 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U13 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U384 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U385 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
assign op_hcompute_conv_stencil_2_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_2_port_controller_flush = flush;
affine_controller__U381 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_2_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_2_port_controller_flush),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U382 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U383 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U386 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U387 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U393_out;
op_hcompute_conv_stencil_3_exe_start_pt__U391 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U402_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U402_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U402_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U402_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U402_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U394 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
assign op_hcompute_conv_stencil_3_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_3_port_controller_flush = flush;
affine_controller__U388 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_3_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_3_port_controller_flush),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U389 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U390 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U426_out;
op_hcompute_conv_stencil_3_write_start_pt__U409 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U540_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U540_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U540_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U540_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U540_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U427 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U68_out;
op_hcompute_conv_stencil_4_exe_start_pt__U66 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U77_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U77_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U77_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U77_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U77_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U69 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
assign op_hcompute_conv_stencil_4_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_4_port_controller_flush = flush;
affine_controller__U63 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_4_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_4_port_controller_flush),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U64 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U65 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U101_out;
op_hcompute_conv_stencil_4_write_start_pt__U84 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U215_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U215_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U215_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U215_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U215_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U102 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U227_out;
op_hcompute_conv_stencil_5_exe_start_pt__U225 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U236_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U236_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U236_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U236_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U236_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U228 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
assign op_hcompute_conv_stencil_5_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_5_port_controller_flush = flush;
affine_controller__U222 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_5_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_5_port_controller_flush),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U223 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U224 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U260_out;
op_hcompute_conv_stencil_5_write_start_pt__U243 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U374_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U374_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U374_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U374_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U374_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U261 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U17 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U18 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
assign op_hcompute_conv_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_conv_stencil_port_controller_flush = flush;
affine_controller__U14 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .rst_n(op_hcompute_conv_stencil_port_controller_rst_n),
    .flush(op_hcompute_conv_stencil_port_controller_flush),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U15 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U16 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U19 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U20 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U3 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U4 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U0 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_input_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_input_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U1 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U2 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U5 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U6 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U59 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U60 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush = flush;
affine_controller__U56 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_flush),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U57 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U58 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U61 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U62 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U26_out;
op_hcompute_hw_output_stencil_exe_start_pt__U24 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U34_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U34_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U34_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U34_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U27 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
assign op_hcompute_hw_output_stencil_port_controller_rst_n = rst_n;
assign op_hcompute_hw_output_stencil_port_controller_flush = flush;
affine_controller__U21 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .rst_n(op_hcompute_hw_output_stencil_port_controller_rst_n),
    .flush(op_hcompute_hw_output_stencil_port_controller_flush),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U22 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U23 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U42_out;
op_hcompute_hw_output_stencil_write_start_pt__U40 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U50_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U50_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U50_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U50_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U43 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

