module inner_sram__U384(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U417(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U450(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U483(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U528(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U601(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U672(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U731(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U791(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
module inner_sram__U832(input logic clk, input logic flush, input logic rst_n, output logic [15:0] rdata, output logic [15:0] wdata, output logic [15:0] raddr, output logic [15:0] waddr, output logic ren_in, output logic wen_in);

  LakeTop lake(.clk(clk), .flush(flush), .rst_n(rst_n), .data_out(rdata), .data_in(wdata), .raddr(raddr), .waddr(waddr), .ren_in(ren_in), .wen_in(wen_in), .clk_en(1), .tile_en(1));

endmodule
