// Module `hw_kernel_global_wrapper_stencil_ub` defined externally
// Module `hw_input_global_wrapper_stencil_ub` defined externally
// Module `conv_stencil_ub` defined externally
module op_hcompute_hw_output_stencil_write_start_pt__U110 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_write_start_control_vars_pt__U113 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_read_start_pt__U92 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_read_start_control_vars_pt__U93 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_output_stencil_exe_start_pt__U94 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U97 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U348 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U349 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U344 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U345 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U346 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U347 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U753 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U754 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U749 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U750 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U751 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U752 (
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_write_start_pt__U21 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_write_start_control_vars_pt__U22 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_read_start_pt__U17 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_read_start_control_vars_pt__U18 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_exe_start_pt__U19 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_exe_start_control_vars_pt__U20 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_write_start_pt__U176 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_write_start_control_vars_pt__U194 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_read_start_pt__U156 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_read_start_control_vars_pt__U157 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_5_exe_start_pt__U158 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U161 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_write_start_pt__U400 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_write_start_control_vars_pt__U418 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_read_start_pt__U380 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_read_start_control_vars_pt__U381 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_4_exe_start_pt__U382 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U385 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_write_start_pt__U588 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_write_start_control_vars_pt__U606 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_read_start_pt__U568 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_read_start_control_vars_pt__U569 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_3_exe_start_pt__U570 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U573 (
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
assign out[4] = in[4];
assign out[3] = in[3];
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_write_start_pt__U67 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_write_start_control_vars_pt__U68 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_read_start_pt__U63 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_read_start_control_vars_pt__U64 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_2_exe_start_pt__U65 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U66 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_write_start_pt__U44 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_write_start_control_vars_pt__U45 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_read_start_pt__U40 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_read_start_control_vars_pt__U41 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module op_hcompute_conv_stencil_1_exe_start_pt__U42 (
    input in,
    output out
);
assign out = in;
endmodule

module op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U43 (
    input [15:0] in [2:0],
    output [15:0] out [2:0]
);
assign out[2] = in[2];
assign out[1] = in[1];
assign out[0] = in[0];
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = in;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    parameter init = 16'h0000
) (
    input [15:0] in,
    input clk,
    output [15:0] out,
    input en
);
wire reg0_clk;
wire [15:0] reg0_in;
assign reg0_clk = clk;
assign reg0_in = en ? in : out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(init),
    .width(16)
) reg0 (
    .clk(reg0_clk),
    .in(reg0_in),
    .out(out)
);
endmodule

module corebit_reg #(
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input in,
    output out
);
reg outReg = init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;
endmodule

module array_delay_U99 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U102_in;
wire _U102_clk;
wire [15:0] _U102_out;
wire [15:0] _U103_in;
wire _U103_clk;
wire [15:0] _U103_out;
assign _U100_in = in[0];
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = in[1];
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U102_in = in[2];
assign _U102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U102_in),
    .clk(_U102_clk),
    .out(_U102_out)
);
assign _U103_in = in[3];
assign _U103_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U103 (
    .in(_U103_in),
    .clk(_U103_clk),
    .out(_U103_out)
);
assign out[3] = _U103_out;
assign out[2] = _U102_out;
assign out[1] = _U101_out;
assign out[0] = _U100_out;
endmodule

module array_delay_U720 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U721_in;
wire _U721_clk;
wire [15:0] _U721_out;
wire [15:0] _U722_in;
wire _U722_clk;
wire [15:0] _U722_out;
wire [15:0] _U723_in;
wire _U723_clk;
wire [15:0] _U723_out;
wire [15:0] _U724_in;
wire _U724_clk;
wire [15:0] _U724_out;
wire [15:0] _U725_in;
wire _U725_clk;
wire [15:0] _U725_out;
assign _U721_in = in[0];
assign _U721_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U721 (
    .in(_U721_in),
    .clk(_U721_clk),
    .out(_U721_out)
);
assign _U722_in = in[1];
assign _U722_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U722 (
    .in(_U722_in),
    .clk(_U722_clk),
    .out(_U722_out)
);
assign _U723_in = in[2];
assign _U723_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U723 (
    .in(_U723_in),
    .clk(_U723_clk),
    .out(_U723_out)
);
assign _U724_in = in[3];
assign _U724_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U724 (
    .in(_U724_in),
    .clk(_U724_clk),
    .out(_U724_out)
);
assign _U725_in = in[4];
assign _U725_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U725 (
    .in(_U725_in),
    .clk(_U725_clk),
    .out(_U725_out)
);
assign out[4] = _U725_out;
assign out[3] = _U724_out;
assign out[2] = _U723_out;
assign out[1] = _U722_out;
assign out[0] = _U721_out;
endmodule

module array_delay_U713 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U714_in;
wire _U714_clk;
wire [15:0] _U714_out;
wire [15:0] _U715_in;
wire _U715_clk;
wire [15:0] _U715_out;
wire [15:0] _U716_in;
wire _U716_clk;
wire [15:0] _U716_out;
wire [15:0] _U717_in;
wire _U717_clk;
wire [15:0] _U717_out;
wire [15:0] _U718_in;
wire _U718_clk;
wire [15:0] _U718_out;
assign _U714_in = in[0];
assign _U714_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U714 (
    .in(_U714_in),
    .clk(_U714_clk),
    .out(_U714_out)
);
assign _U715_in = in[1];
assign _U715_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U715 (
    .in(_U715_in),
    .clk(_U715_clk),
    .out(_U715_out)
);
assign _U716_in = in[2];
assign _U716_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U716 (
    .in(_U716_in),
    .clk(_U716_clk),
    .out(_U716_out)
);
assign _U717_in = in[3];
assign _U717_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U717 (
    .in(_U717_in),
    .clk(_U717_clk),
    .out(_U717_out)
);
assign _U718_in = in[4];
assign _U718_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U718 (
    .in(_U718_in),
    .clk(_U718_clk),
    .out(_U718_out)
);
assign out[4] = _U718_out;
assign out[3] = _U717_out;
assign out[2] = _U716_out;
assign out[1] = _U715_out;
assign out[0] = _U714_out;
endmodule

module array_delay_U706 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U707_in;
wire _U707_clk;
wire [15:0] _U707_out;
wire [15:0] _U708_in;
wire _U708_clk;
wire [15:0] _U708_out;
wire [15:0] _U709_in;
wire _U709_clk;
wire [15:0] _U709_out;
wire [15:0] _U710_in;
wire _U710_clk;
wire [15:0] _U710_out;
wire [15:0] _U711_in;
wire _U711_clk;
wire [15:0] _U711_out;
assign _U707_in = in[0];
assign _U707_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U707 (
    .in(_U707_in),
    .clk(_U707_clk),
    .out(_U707_out)
);
assign _U708_in = in[1];
assign _U708_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U708 (
    .in(_U708_in),
    .clk(_U708_clk),
    .out(_U708_out)
);
assign _U709_in = in[2];
assign _U709_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U709 (
    .in(_U709_in),
    .clk(_U709_clk),
    .out(_U709_out)
);
assign _U710_in = in[3];
assign _U710_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U710 (
    .in(_U710_in),
    .clk(_U710_clk),
    .out(_U710_out)
);
assign _U711_in = in[4];
assign _U711_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U711 (
    .in(_U711_in),
    .clk(_U711_clk),
    .out(_U711_out)
);
assign out[4] = _U711_out;
assign out[3] = _U710_out;
assign out[2] = _U709_out;
assign out[1] = _U708_out;
assign out[0] = _U707_out;
endmodule

module array_delay_U699 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U700_in;
wire _U700_clk;
wire [15:0] _U700_out;
wire [15:0] _U701_in;
wire _U701_clk;
wire [15:0] _U701_out;
wire [15:0] _U702_in;
wire _U702_clk;
wire [15:0] _U702_out;
wire [15:0] _U703_in;
wire _U703_clk;
wire [15:0] _U703_out;
wire [15:0] _U704_in;
wire _U704_clk;
wire [15:0] _U704_out;
assign _U700_in = in[0];
assign _U700_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U700 (
    .in(_U700_in),
    .clk(_U700_clk),
    .out(_U700_out)
);
assign _U701_in = in[1];
assign _U701_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U701 (
    .in(_U701_in),
    .clk(_U701_clk),
    .out(_U701_out)
);
assign _U702_in = in[2];
assign _U702_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U702 (
    .in(_U702_in),
    .clk(_U702_clk),
    .out(_U702_out)
);
assign _U703_in = in[3];
assign _U703_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U703 (
    .in(_U703_in),
    .clk(_U703_clk),
    .out(_U703_out)
);
assign _U704_in = in[4];
assign _U704_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U704 (
    .in(_U704_in),
    .clk(_U704_clk),
    .out(_U704_out)
);
assign out[4] = _U704_out;
assign out[3] = _U703_out;
assign out[2] = _U702_out;
assign out[1] = _U701_out;
assign out[0] = _U700_out;
endmodule

module array_delay_U692 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U693_in;
wire _U693_clk;
wire [15:0] _U693_out;
wire [15:0] _U694_in;
wire _U694_clk;
wire [15:0] _U694_out;
wire [15:0] _U695_in;
wire _U695_clk;
wire [15:0] _U695_out;
wire [15:0] _U696_in;
wire _U696_clk;
wire [15:0] _U696_out;
wire [15:0] _U697_in;
wire _U697_clk;
wire [15:0] _U697_out;
assign _U693_in = in[0];
assign _U693_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U693 (
    .in(_U693_in),
    .clk(_U693_clk),
    .out(_U693_out)
);
assign _U694_in = in[1];
assign _U694_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U694 (
    .in(_U694_in),
    .clk(_U694_clk),
    .out(_U694_out)
);
assign _U695_in = in[2];
assign _U695_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U695 (
    .in(_U695_in),
    .clk(_U695_clk),
    .out(_U695_out)
);
assign _U696_in = in[3];
assign _U696_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U696 (
    .in(_U696_in),
    .clk(_U696_clk),
    .out(_U696_out)
);
assign _U697_in = in[4];
assign _U697_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U697 (
    .in(_U697_in),
    .clk(_U697_clk),
    .out(_U697_out)
);
assign out[4] = _U697_out;
assign out[3] = _U696_out;
assign out[2] = _U695_out;
assign out[1] = _U694_out;
assign out[0] = _U693_out;
endmodule

module array_delay_U685 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U686_in;
wire _U686_clk;
wire [15:0] _U686_out;
wire [15:0] _U687_in;
wire _U687_clk;
wire [15:0] _U687_out;
wire [15:0] _U688_in;
wire _U688_clk;
wire [15:0] _U688_out;
wire [15:0] _U689_in;
wire _U689_clk;
wire [15:0] _U689_out;
wire [15:0] _U690_in;
wire _U690_clk;
wire [15:0] _U690_out;
assign _U686_in = in[0];
assign _U686_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U686 (
    .in(_U686_in),
    .clk(_U686_clk),
    .out(_U686_out)
);
assign _U687_in = in[1];
assign _U687_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U687 (
    .in(_U687_in),
    .clk(_U687_clk),
    .out(_U687_out)
);
assign _U688_in = in[2];
assign _U688_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U688 (
    .in(_U688_in),
    .clk(_U688_clk),
    .out(_U688_out)
);
assign _U689_in = in[3];
assign _U689_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U689 (
    .in(_U689_in),
    .clk(_U689_clk),
    .out(_U689_out)
);
assign _U690_in = in[4];
assign _U690_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U690 (
    .in(_U690_in),
    .clk(_U690_clk),
    .out(_U690_out)
);
assign out[4] = _U690_out;
assign out[3] = _U689_out;
assign out[2] = _U688_out;
assign out[1] = _U687_out;
assign out[0] = _U686_out;
endmodule

module array_delay_U678 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U679_in;
wire _U679_clk;
wire [15:0] _U679_out;
wire [15:0] _U680_in;
wire _U680_clk;
wire [15:0] _U680_out;
wire [15:0] _U681_in;
wire _U681_clk;
wire [15:0] _U681_out;
wire [15:0] _U682_in;
wire _U682_clk;
wire [15:0] _U682_out;
wire [15:0] _U683_in;
wire _U683_clk;
wire [15:0] _U683_out;
assign _U679_in = in[0];
assign _U679_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U679 (
    .in(_U679_in),
    .clk(_U679_clk),
    .out(_U679_out)
);
assign _U680_in = in[1];
assign _U680_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U680 (
    .in(_U680_in),
    .clk(_U680_clk),
    .out(_U680_out)
);
assign _U681_in = in[2];
assign _U681_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U681 (
    .in(_U681_in),
    .clk(_U681_clk),
    .out(_U681_out)
);
assign _U682_in = in[3];
assign _U682_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U682 (
    .in(_U682_in),
    .clk(_U682_clk),
    .out(_U682_out)
);
assign _U683_in = in[4];
assign _U683_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U683 (
    .in(_U683_in),
    .clk(_U683_clk),
    .out(_U683_out)
);
assign out[4] = _U683_out;
assign out[3] = _U682_out;
assign out[2] = _U681_out;
assign out[1] = _U680_out;
assign out[0] = _U679_out;
endmodule

module array_delay_U671 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U672_in;
wire _U672_clk;
wire [15:0] _U672_out;
wire [15:0] _U673_in;
wire _U673_clk;
wire [15:0] _U673_out;
wire [15:0] _U674_in;
wire _U674_clk;
wire [15:0] _U674_out;
wire [15:0] _U675_in;
wire _U675_clk;
wire [15:0] _U675_out;
wire [15:0] _U676_in;
wire _U676_clk;
wire [15:0] _U676_out;
assign _U672_in = in[0];
assign _U672_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U672 (
    .in(_U672_in),
    .clk(_U672_clk),
    .out(_U672_out)
);
assign _U673_in = in[1];
assign _U673_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U673 (
    .in(_U673_in),
    .clk(_U673_clk),
    .out(_U673_out)
);
assign _U674_in = in[2];
assign _U674_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U674 (
    .in(_U674_in),
    .clk(_U674_clk),
    .out(_U674_out)
);
assign _U675_in = in[3];
assign _U675_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U675 (
    .in(_U675_in),
    .clk(_U675_clk),
    .out(_U675_out)
);
assign _U676_in = in[4];
assign _U676_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U676 (
    .in(_U676_in),
    .clk(_U676_clk),
    .out(_U676_out)
);
assign out[4] = _U676_out;
assign out[3] = _U675_out;
assign out[2] = _U674_out;
assign out[1] = _U673_out;
assign out[0] = _U672_out;
endmodule

module array_delay_U664 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U665_in;
wire _U665_clk;
wire [15:0] _U665_out;
wire [15:0] _U666_in;
wire _U666_clk;
wire [15:0] _U666_out;
wire [15:0] _U667_in;
wire _U667_clk;
wire [15:0] _U667_out;
wire [15:0] _U668_in;
wire _U668_clk;
wire [15:0] _U668_out;
wire [15:0] _U669_in;
wire _U669_clk;
wire [15:0] _U669_out;
assign _U665_in = in[0];
assign _U665_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U665 (
    .in(_U665_in),
    .clk(_U665_clk),
    .out(_U665_out)
);
assign _U666_in = in[1];
assign _U666_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U666 (
    .in(_U666_in),
    .clk(_U666_clk),
    .out(_U666_out)
);
assign _U667_in = in[2];
assign _U667_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U667 (
    .in(_U667_in),
    .clk(_U667_clk),
    .out(_U667_out)
);
assign _U668_in = in[3];
assign _U668_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U668 (
    .in(_U668_in),
    .clk(_U668_clk),
    .out(_U668_out)
);
assign _U669_in = in[4];
assign _U669_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U669 (
    .in(_U669_in),
    .clk(_U669_clk),
    .out(_U669_out)
);
assign out[4] = _U669_out;
assign out[3] = _U668_out;
assign out[2] = _U667_out;
assign out[1] = _U666_out;
assign out[0] = _U665_out;
endmodule

module array_delay_U657 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U658_in;
wire _U658_clk;
wire [15:0] _U658_out;
wire [15:0] _U659_in;
wire _U659_clk;
wire [15:0] _U659_out;
wire [15:0] _U660_in;
wire _U660_clk;
wire [15:0] _U660_out;
wire [15:0] _U661_in;
wire _U661_clk;
wire [15:0] _U661_out;
wire [15:0] _U662_in;
wire _U662_clk;
wire [15:0] _U662_out;
assign _U658_in = in[0];
assign _U658_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U658 (
    .in(_U658_in),
    .clk(_U658_clk),
    .out(_U658_out)
);
assign _U659_in = in[1];
assign _U659_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U659 (
    .in(_U659_in),
    .clk(_U659_clk),
    .out(_U659_out)
);
assign _U660_in = in[2];
assign _U660_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U660 (
    .in(_U660_in),
    .clk(_U660_clk),
    .out(_U660_out)
);
assign _U661_in = in[3];
assign _U661_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U661 (
    .in(_U661_in),
    .clk(_U661_clk),
    .out(_U661_out)
);
assign _U662_in = in[4];
assign _U662_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U662 (
    .in(_U662_in),
    .clk(_U662_clk),
    .out(_U662_out)
);
assign out[4] = _U662_out;
assign out[3] = _U661_out;
assign out[2] = _U660_out;
assign out[1] = _U659_out;
assign out[0] = _U658_out;
endmodule

module array_delay_U650 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U651_in;
wire _U651_clk;
wire [15:0] _U651_out;
wire [15:0] _U652_in;
wire _U652_clk;
wire [15:0] _U652_out;
wire [15:0] _U653_in;
wire _U653_clk;
wire [15:0] _U653_out;
wire [15:0] _U654_in;
wire _U654_clk;
wire [15:0] _U654_out;
wire [15:0] _U655_in;
wire _U655_clk;
wire [15:0] _U655_out;
assign _U651_in = in[0];
assign _U651_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U651 (
    .in(_U651_in),
    .clk(_U651_clk),
    .out(_U651_out)
);
assign _U652_in = in[1];
assign _U652_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U652 (
    .in(_U652_in),
    .clk(_U652_clk),
    .out(_U652_out)
);
assign _U653_in = in[2];
assign _U653_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U653 (
    .in(_U653_in),
    .clk(_U653_clk),
    .out(_U653_out)
);
assign _U654_in = in[3];
assign _U654_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U654 (
    .in(_U654_in),
    .clk(_U654_clk),
    .out(_U654_out)
);
assign _U655_in = in[4];
assign _U655_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U655 (
    .in(_U655_in),
    .clk(_U655_clk),
    .out(_U655_out)
);
assign out[4] = _U655_out;
assign out[3] = _U654_out;
assign out[2] = _U653_out;
assign out[1] = _U652_out;
assign out[0] = _U651_out;
endmodule

module array_delay_U643 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U644_in;
wire _U644_clk;
wire [15:0] _U644_out;
wire [15:0] _U645_in;
wire _U645_clk;
wire [15:0] _U645_out;
wire [15:0] _U646_in;
wire _U646_clk;
wire [15:0] _U646_out;
wire [15:0] _U647_in;
wire _U647_clk;
wire [15:0] _U647_out;
wire [15:0] _U648_in;
wire _U648_clk;
wire [15:0] _U648_out;
assign _U644_in = in[0];
assign _U644_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U644 (
    .in(_U644_in),
    .clk(_U644_clk),
    .out(_U644_out)
);
assign _U645_in = in[1];
assign _U645_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U645 (
    .in(_U645_in),
    .clk(_U645_clk),
    .out(_U645_out)
);
assign _U646_in = in[2];
assign _U646_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U646 (
    .in(_U646_in),
    .clk(_U646_clk),
    .out(_U646_out)
);
assign _U647_in = in[3];
assign _U647_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U647 (
    .in(_U647_in),
    .clk(_U647_clk),
    .out(_U647_out)
);
assign _U648_in = in[4];
assign _U648_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U648 (
    .in(_U648_in),
    .clk(_U648_clk),
    .out(_U648_out)
);
assign out[4] = _U648_out;
assign out[3] = _U647_out;
assign out[2] = _U646_out;
assign out[1] = _U645_out;
assign out[0] = _U644_out;
endmodule

module array_delay_U636 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U637_in;
wire _U637_clk;
wire [15:0] _U637_out;
wire [15:0] _U638_in;
wire _U638_clk;
wire [15:0] _U638_out;
wire [15:0] _U639_in;
wire _U639_clk;
wire [15:0] _U639_out;
wire [15:0] _U640_in;
wire _U640_clk;
wire [15:0] _U640_out;
wire [15:0] _U641_in;
wire _U641_clk;
wire [15:0] _U641_out;
assign _U637_in = in[0];
assign _U637_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U637 (
    .in(_U637_in),
    .clk(_U637_clk),
    .out(_U637_out)
);
assign _U638_in = in[1];
assign _U638_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U638 (
    .in(_U638_in),
    .clk(_U638_clk),
    .out(_U638_out)
);
assign _U639_in = in[2];
assign _U639_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U639 (
    .in(_U639_in),
    .clk(_U639_clk),
    .out(_U639_out)
);
assign _U640_in = in[3];
assign _U640_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U640 (
    .in(_U640_in),
    .clk(_U640_clk),
    .out(_U640_out)
);
assign _U641_in = in[4];
assign _U641_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U641 (
    .in(_U641_in),
    .clk(_U641_clk),
    .out(_U641_out)
);
assign out[4] = _U641_out;
assign out[3] = _U640_out;
assign out[2] = _U639_out;
assign out[1] = _U638_out;
assign out[0] = _U637_out;
endmodule

module array_delay_U629 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U630_in;
wire _U630_clk;
wire [15:0] _U630_out;
wire [15:0] _U631_in;
wire _U631_clk;
wire [15:0] _U631_out;
wire [15:0] _U632_in;
wire _U632_clk;
wire [15:0] _U632_out;
wire [15:0] _U633_in;
wire _U633_clk;
wire [15:0] _U633_out;
wire [15:0] _U634_in;
wire _U634_clk;
wire [15:0] _U634_out;
assign _U630_in = in[0];
assign _U630_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U630 (
    .in(_U630_in),
    .clk(_U630_clk),
    .out(_U630_out)
);
assign _U631_in = in[1];
assign _U631_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U631 (
    .in(_U631_in),
    .clk(_U631_clk),
    .out(_U631_out)
);
assign _U632_in = in[2];
assign _U632_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U632 (
    .in(_U632_in),
    .clk(_U632_clk),
    .out(_U632_out)
);
assign _U633_in = in[3];
assign _U633_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U633 (
    .in(_U633_in),
    .clk(_U633_clk),
    .out(_U633_out)
);
assign _U634_in = in[4];
assign _U634_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U634 (
    .in(_U634_in),
    .clk(_U634_clk),
    .out(_U634_out)
);
assign out[4] = _U634_out;
assign out[3] = _U633_out;
assign out[2] = _U632_out;
assign out[1] = _U631_out;
assign out[0] = _U630_out;
endmodule

module array_delay_U622 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U623_in;
wire _U623_clk;
wire [15:0] _U623_out;
wire [15:0] _U624_in;
wire _U624_clk;
wire [15:0] _U624_out;
wire [15:0] _U625_in;
wire _U625_clk;
wire [15:0] _U625_out;
wire [15:0] _U626_in;
wire _U626_clk;
wire [15:0] _U626_out;
wire [15:0] _U627_in;
wire _U627_clk;
wire [15:0] _U627_out;
assign _U623_in = in[0];
assign _U623_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U623 (
    .in(_U623_in),
    .clk(_U623_clk),
    .out(_U623_out)
);
assign _U624_in = in[1];
assign _U624_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U624 (
    .in(_U624_in),
    .clk(_U624_clk),
    .out(_U624_out)
);
assign _U625_in = in[2];
assign _U625_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U625 (
    .in(_U625_in),
    .clk(_U625_clk),
    .out(_U625_out)
);
assign _U626_in = in[3];
assign _U626_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U626 (
    .in(_U626_in),
    .clk(_U626_clk),
    .out(_U626_out)
);
assign _U627_in = in[4];
assign _U627_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U627 (
    .in(_U627_in),
    .clk(_U627_clk),
    .out(_U627_out)
);
assign out[4] = _U627_out;
assign out[3] = _U626_out;
assign out[2] = _U625_out;
assign out[1] = _U624_out;
assign out[0] = _U623_out;
endmodule

module array_delay_U615 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U616_in;
wire _U616_clk;
wire [15:0] _U616_out;
wire [15:0] _U617_in;
wire _U617_clk;
wire [15:0] _U617_out;
wire [15:0] _U618_in;
wire _U618_clk;
wire [15:0] _U618_out;
wire [15:0] _U619_in;
wire _U619_clk;
wire [15:0] _U619_out;
wire [15:0] _U620_in;
wire _U620_clk;
wire [15:0] _U620_out;
assign _U616_in = in[0];
assign _U616_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U616 (
    .in(_U616_in),
    .clk(_U616_clk),
    .out(_U616_out)
);
assign _U617_in = in[1];
assign _U617_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U617 (
    .in(_U617_in),
    .clk(_U617_clk),
    .out(_U617_out)
);
assign _U618_in = in[2];
assign _U618_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U618 (
    .in(_U618_in),
    .clk(_U618_clk),
    .out(_U618_out)
);
assign _U619_in = in[3];
assign _U619_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U619 (
    .in(_U619_in),
    .clk(_U619_clk),
    .out(_U619_out)
);
assign _U620_in = in[4];
assign _U620_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U620 (
    .in(_U620_in),
    .clk(_U620_clk),
    .out(_U620_out)
);
assign out[4] = _U620_out;
assign out[3] = _U619_out;
assign out[2] = _U618_out;
assign out[1] = _U617_out;
assign out[0] = _U616_out;
endmodule

module array_delay_U608 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
wire [15:0] _U611_in;
wire _U611_clk;
wire [15:0] _U611_out;
wire [15:0] _U612_in;
wire _U612_clk;
wire [15:0] _U612_out;
wire [15:0] _U613_in;
wire _U613_clk;
wire [15:0] _U613_out;
assign _U609_in = in[0];
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = in[1];
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
assign _U611_in = in[2];
assign _U611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U611 (
    .in(_U611_in),
    .clk(_U611_clk),
    .out(_U611_out)
);
assign _U612_in = in[3];
assign _U612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U612 (
    .in(_U612_in),
    .clk(_U612_clk),
    .out(_U612_out)
);
assign _U613_in = in[4];
assign _U613_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U613 (
    .in(_U613_in),
    .clk(_U613_clk),
    .out(_U613_out)
);
assign out[4] = _U613_out;
assign out[3] = _U612_out;
assign out[2] = _U611_out;
assign out[1] = _U610_out;
assign out[0] = _U609_out;
endmodule

module array_delay_U582 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
wire [15:0] _U585_in;
wire _U585_clk;
wire [15:0] _U585_out;
wire [15:0] _U586_in;
wire _U586_clk;
wire [15:0] _U586_out;
wire [15:0] _U587_in;
wire _U587_clk;
wire [15:0] _U587_out;
assign _U583_in = in[0];
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = in[1];
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign _U585_in = in[2];
assign _U585_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U585 (
    .in(_U585_in),
    .clk(_U585_clk),
    .out(_U585_out)
);
assign _U586_in = in[3];
assign _U586_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U586 (
    .in(_U586_in),
    .clk(_U586_clk),
    .out(_U586_out)
);
assign _U587_in = in[4];
assign _U587_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U587 (
    .in(_U587_in),
    .clk(_U587_clk),
    .out(_U587_out)
);
assign out[4] = _U587_out;
assign out[3] = _U586_out;
assign out[2] = _U585_out;
assign out[1] = _U584_out;
assign out[0] = _U583_out;
endmodule

module array_delay_U575 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U576_in;
wire _U576_clk;
wire [15:0] _U576_out;
wire [15:0] _U577_in;
wire _U577_clk;
wire [15:0] _U577_out;
wire [15:0] _U578_in;
wire _U578_clk;
wire [15:0] _U578_out;
wire [15:0] _U579_in;
wire _U579_clk;
wire [15:0] _U579_out;
wire [15:0] _U580_in;
wire _U580_clk;
wire [15:0] _U580_out;
assign _U576_in = in[0];
assign _U576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U576_in),
    .clk(_U576_clk),
    .out(_U576_out)
);
assign _U577_in = in[1];
assign _U577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U577 (
    .in(_U577_in),
    .clk(_U577_clk),
    .out(_U577_out)
);
assign _U578_in = in[2];
assign _U578_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U578 (
    .in(_U578_in),
    .clk(_U578_clk),
    .out(_U578_out)
);
assign _U579_in = in[3];
assign _U579_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U579 (
    .in(_U579_in),
    .clk(_U579_clk),
    .out(_U579_out)
);
assign _U580_in = in[4];
assign _U580_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U580 (
    .in(_U580_in),
    .clk(_U580_clk),
    .out(_U580_out)
);
assign out[4] = _U580_out;
assign out[3] = _U579_out;
assign out[2] = _U578_out;
assign out[1] = _U577_out;
assign out[0] = _U576_out;
endmodule

module array_delay_U532 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U533_in;
wire _U533_clk;
wire [15:0] _U533_out;
wire [15:0] _U534_in;
wire _U534_clk;
wire [15:0] _U534_out;
wire [15:0] _U535_in;
wire _U535_clk;
wire [15:0] _U535_out;
wire [15:0] _U536_in;
wire _U536_clk;
wire [15:0] _U536_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
assign _U533_in = in[0];
assign _U533_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U533 (
    .in(_U533_in),
    .clk(_U533_clk),
    .out(_U533_out)
);
assign _U534_in = in[1];
assign _U534_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U534 (
    .in(_U534_in),
    .clk(_U534_clk),
    .out(_U534_out)
);
assign _U535_in = in[2];
assign _U535_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U535 (
    .in(_U535_in),
    .clk(_U535_clk),
    .out(_U535_out)
);
assign _U536_in = in[3];
assign _U536_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U536 (
    .in(_U536_in),
    .clk(_U536_clk),
    .out(_U536_out)
);
assign _U537_in = in[4];
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign out[4] = _U537_out;
assign out[3] = _U536_out;
assign out[2] = _U535_out;
assign out[1] = _U534_out;
assign out[0] = _U533_out;
endmodule

module array_delay_U525 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U526_in;
wire _U526_clk;
wire [15:0] _U526_out;
wire [15:0] _U527_in;
wire _U527_clk;
wire [15:0] _U527_out;
wire [15:0] _U528_in;
wire _U528_clk;
wire [15:0] _U528_out;
wire [15:0] _U529_in;
wire _U529_clk;
wire [15:0] _U529_out;
wire [15:0] _U530_in;
wire _U530_clk;
wire [15:0] _U530_out;
assign _U526_in = in[0];
assign _U526_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U526 (
    .in(_U526_in),
    .clk(_U526_clk),
    .out(_U526_out)
);
assign _U527_in = in[1];
assign _U527_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U527 (
    .in(_U527_in),
    .clk(_U527_clk),
    .out(_U527_out)
);
assign _U528_in = in[2];
assign _U528_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U528 (
    .in(_U528_in),
    .clk(_U528_clk),
    .out(_U528_out)
);
assign _U529_in = in[3];
assign _U529_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U529 (
    .in(_U529_in),
    .clk(_U529_clk),
    .out(_U529_out)
);
assign _U530_in = in[4];
assign _U530_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U530 (
    .in(_U530_in),
    .clk(_U530_clk),
    .out(_U530_out)
);
assign out[4] = _U530_out;
assign out[3] = _U529_out;
assign out[2] = _U528_out;
assign out[1] = _U527_out;
assign out[0] = _U526_out;
endmodule

module array_delay_U518 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire _U520_clk;
wire [15:0] _U520_out;
wire [15:0] _U521_in;
wire _U521_clk;
wire [15:0] _U521_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
assign _U519_in = in[0];
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = in[1];
assign _U520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U520_in),
    .clk(_U520_clk),
    .out(_U520_out)
);
assign _U521_in = in[2];
assign _U521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U521_in),
    .clk(_U521_clk),
    .out(_U521_out)
);
assign _U522_in = in[3];
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = in[4];
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign out[4] = _U523_out;
assign out[3] = _U522_out;
assign out[2] = _U521_out;
assign out[1] = _U520_out;
assign out[0] = _U519_out;
endmodule

module array_delay_U511 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire _U513_clk;
wire [15:0] _U513_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
assign _U512_in = in[0];
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = in[1];
assign _U513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U513_in),
    .clk(_U513_clk),
    .out(_U513_out)
);
assign _U514_in = in[2];
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = in[3];
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = in[4];
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign out[4] = _U516_out;
assign out[3] = _U515_out;
assign out[2] = _U514_out;
assign out[1] = _U513_out;
assign out[0] = _U512_out;
endmodule

module array_delay_U504 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire _U506_clk;
wire [15:0] _U506_out;
wire [15:0] _U507_in;
wire _U507_clk;
wire [15:0] _U507_out;
wire [15:0] _U508_in;
wire _U508_clk;
wire [15:0] _U508_out;
wire [15:0] _U509_in;
wire _U509_clk;
wire [15:0] _U509_out;
assign _U505_in = in[0];
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = in[1];
assign _U506_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U506 (
    .in(_U506_in),
    .clk(_U506_clk),
    .out(_U506_out)
);
assign _U507_in = in[2];
assign _U507_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U507 (
    .in(_U507_in),
    .clk(_U507_clk),
    .out(_U507_out)
);
assign _U508_in = in[3];
assign _U508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U508 (
    .in(_U508_in),
    .clk(_U508_clk),
    .out(_U508_out)
);
assign _U509_in = in[4];
assign _U509_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U509 (
    .in(_U509_in),
    .clk(_U509_clk),
    .out(_U509_out)
);
assign out[4] = _U509_out;
assign out[3] = _U508_out;
assign out[2] = _U507_out;
assign out[1] = _U506_out;
assign out[0] = _U505_out;
endmodule

module array_delay_U497 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U498_in;
wire _U498_clk;
wire [15:0] _U498_out;
wire [15:0] _U499_in;
wire _U499_clk;
wire [15:0] _U499_out;
wire [15:0] _U500_in;
wire _U500_clk;
wire [15:0] _U500_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire _U502_clk;
wire [15:0] _U502_out;
assign _U498_in = in[0];
assign _U498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U498_in),
    .clk(_U498_clk),
    .out(_U498_out)
);
assign _U499_in = in[1];
assign _U499_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U499 (
    .in(_U499_in),
    .clk(_U499_clk),
    .out(_U499_out)
);
assign _U500_in = in[2];
assign _U500_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U500 (
    .in(_U500_in),
    .clk(_U500_clk),
    .out(_U500_out)
);
assign _U501_in = in[3];
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = in[4];
assign _U502_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U502 (
    .in(_U502_in),
    .clk(_U502_clk),
    .out(_U502_out)
);
assign out[4] = _U502_out;
assign out[3] = _U501_out;
assign out[2] = _U500_out;
assign out[1] = _U499_out;
assign out[0] = _U498_out;
endmodule

module array_delay_U490 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U491_in;
wire _U491_clk;
wire [15:0] _U491_out;
wire [15:0] _U492_in;
wire _U492_clk;
wire [15:0] _U492_out;
wire [15:0] _U493_in;
wire _U493_clk;
wire [15:0] _U493_out;
wire [15:0] _U494_in;
wire _U494_clk;
wire [15:0] _U494_out;
wire [15:0] _U495_in;
wire _U495_clk;
wire [15:0] _U495_out;
assign _U491_in = in[0];
assign _U491_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U491 (
    .in(_U491_in),
    .clk(_U491_clk),
    .out(_U491_out)
);
assign _U492_in = in[1];
assign _U492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(_U492_in),
    .clk(_U492_clk),
    .out(_U492_out)
);
assign _U493_in = in[2];
assign _U493_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U493 (
    .in(_U493_in),
    .clk(_U493_clk),
    .out(_U493_out)
);
assign _U494_in = in[3];
assign _U494_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U494 (
    .in(_U494_in),
    .clk(_U494_clk),
    .out(_U494_out)
);
assign _U495_in = in[4];
assign _U495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U495 (
    .in(_U495_in),
    .clk(_U495_clk),
    .out(_U495_out)
);
assign out[4] = _U495_out;
assign out[3] = _U494_out;
assign out[2] = _U493_out;
assign out[1] = _U492_out;
assign out[0] = _U491_out;
endmodule

module array_delay_U483 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U484_in;
wire _U484_clk;
wire [15:0] _U484_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire _U487_clk;
wire [15:0] _U487_out;
wire [15:0] _U488_in;
wire _U488_clk;
wire [15:0] _U488_out;
assign _U484_in = in[0];
assign _U484_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(_U484_in),
    .clk(_U484_clk),
    .out(_U484_out)
);
assign _U485_in = in[1];
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = in[2];
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = in[3];
assign _U487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U487 (
    .in(_U487_in),
    .clk(_U487_clk),
    .out(_U487_out)
);
assign _U488_in = in[4];
assign _U488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U488 (
    .in(_U488_in),
    .clk(_U488_clk),
    .out(_U488_out)
);
assign out[4] = _U488_out;
assign out[3] = _U487_out;
assign out[2] = _U486_out;
assign out[1] = _U485_out;
assign out[0] = _U484_out;
endmodule

module array_delay_U476 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire _U478_clk;
wire [15:0] _U478_out;
wire [15:0] _U479_in;
wire _U479_clk;
wire [15:0] _U479_out;
wire [15:0] _U480_in;
wire _U480_clk;
wire [15:0] _U480_out;
wire [15:0] _U481_in;
wire _U481_clk;
wire [15:0] _U481_out;
assign _U477_in = in[0];
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = in[1];
assign _U478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(_U478_in),
    .clk(_U478_clk),
    .out(_U478_out)
);
assign _U479_in = in[2];
assign _U479_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U479 (
    .in(_U479_in),
    .clk(_U479_clk),
    .out(_U479_out)
);
assign _U480_in = in[3];
assign _U480_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U480 (
    .in(_U480_in),
    .clk(_U480_clk),
    .out(_U480_out)
);
assign _U481_in = in[4];
assign _U481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U481_in),
    .clk(_U481_clk),
    .out(_U481_out)
);
assign out[4] = _U481_out;
assign out[3] = _U480_out;
assign out[2] = _U479_out;
assign out[1] = _U478_out;
assign out[0] = _U477_out;
endmodule

module array_delay_U469 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U470_in;
wire _U470_clk;
wire [15:0] _U470_out;
wire [15:0] _U471_in;
wire _U471_clk;
wire [15:0] _U471_out;
wire [15:0] _U472_in;
wire _U472_clk;
wire [15:0] _U472_out;
wire [15:0] _U473_in;
wire _U473_clk;
wire [15:0] _U473_out;
wire [15:0] _U474_in;
wire _U474_clk;
wire [15:0] _U474_out;
assign _U470_in = in[0];
assign _U470_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U470 (
    .in(_U470_in),
    .clk(_U470_clk),
    .out(_U470_out)
);
assign _U471_in = in[1];
assign _U471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U471 (
    .in(_U471_in),
    .clk(_U471_clk),
    .out(_U471_out)
);
assign _U472_in = in[2];
assign _U472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U472 (
    .in(_U472_in),
    .clk(_U472_clk),
    .out(_U472_out)
);
assign _U473_in = in[3];
assign _U473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U473 (
    .in(_U473_in),
    .clk(_U473_clk),
    .out(_U473_out)
);
assign _U474_in = in[4];
assign _U474_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U474 (
    .in(_U474_in),
    .clk(_U474_clk),
    .out(_U474_out)
);
assign out[4] = _U474_out;
assign out[3] = _U473_out;
assign out[2] = _U472_out;
assign out[1] = _U471_out;
assign out[0] = _U470_out;
endmodule

module array_delay_U462 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U463_in;
wire _U463_clk;
wire [15:0] _U463_out;
wire [15:0] _U464_in;
wire _U464_clk;
wire [15:0] _U464_out;
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire _U466_clk;
wire [15:0] _U466_out;
wire [15:0] _U467_in;
wire _U467_clk;
wire [15:0] _U467_out;
assign _U463_in = in[0];
assign _U463_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U463 (
    .in(_U463_in),
    .clk(_U463_clk),
    .out(_U463_out)
);
assign _U464_in = in[1];
assign _U464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U464 (
    .in(_U464_in),
    .clk(_U464_clk),
    .out(_U464_out)
);
assign _U465_in = in[2];
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = in[3];
assign _U466_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U466 (
    .in(_U466_in),
    .clk(_U466_clk),
    .out(_U466_out)
);
assign _U467_in = in[4];
assign _U467_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U467 (
    .in(_U467_in),
    .clk(_U467_clk),
    .out(_U467_out)
);
assign out[4] = _U467_out;
assign out[3] = _U466_out;
assign out[2] = _U465_out;
assign out[1] = _U464_out;
assign out[0] = _U463_out;
endmodule

module array_delay_U455 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U456_in;
wire _U456_clk;
wire [15:0] _U456_out;
wire [15:0] _U457_in;
wire _U457_clk;
wire [15:0] _U457_out;
wire [15:0] _U458_in;
wire _U458_clk;
wire [15:0] _U458_out;
wire [15:0] _U459_in;
wire _U459_clk;
wire [15:0] _U459_out;
wire [15:0] _U460_in;
wire _U460_clk;
wire [15:0] _U460_out;
assign _U456_in = in[0];
assign _U456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U456 (
    .in(_U456_in),
    .clk(_U456_clk),
    .out(_U456_out)
);
assign _U457_in = in[1];
assign _U457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U457 (
    .in(_U457_in),
    .clk(_U457_clk),
    .out(_U457_out)
);
assign _U458_in = in[2];
assign _U458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U458 (
    .in(_U458_in),
    .clk(_U458_clk),
    .out(_U458_out)
);
assign _U459_in = in[3];
assign _U459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U459 (
    .in(_U459_in),
    .clk(_U459_clk),
    .out(_U459_out)
);
assign _U460_in = in[4];
assign _U460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U460 (
    .in(_U460_in),
    .clk(_U460_clk),
    .out(_U460_out)
);
assign out[4] = _U460_out;
assign out[3] = _U459_out;
assign out[2] = _U458_out;
assign out[1] = _U457_out;
assign out[0] = _U456_out;
endmodule

module array_delay_U448 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U449_in;
wire _U449_clk;
wire [15:0] _U449_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
wire [15:0] _U451_in;
wire _U451_clk;
wire [15:0] _U451_out;
wire [15:0] _U452_in;
wire _U452_clk;
wire [15:0] _U452_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
assign _U449_in = in[0];
assign _U449_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U449 (
    .in(_U449_in),
    .clk(_U449_clk),
    .out(_U449_out)
);
assign _U450_in = in[1];
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign _U451_in = in[2];
assign _U451_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U451 (
    .in(_U451_in),
    .clk(_U451_clk),
    .out(_U451_out)
);
assign _U452_in = in[3];
assign _U452_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U452 (
    .in(_U452_in),
    .clk(_U452_clk),
    .out(_U452_out)
);
assign _U453_in = in[4];
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign out[4] = _U453_out;
assign out[3] = _U452_out;
assign out[2] = _U451_out;
assign out[1] = _U450_out;
assign out[0] = _U449_out;
endmodule

module array_delay_U441 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
assign _U442_in = in[0];
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = in[1];
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = in[2];
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = in[3];
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = in[4];
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign out[4] = _U446_out;
assign out[3] = _U445_out;
assign out[2] = _U444_out;
assign out[1] = _U443_out;
assign out[0] = _U442_out;
endmodule

module array_delay_U434 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U435_in;
wire _U435_clk;
wire [15:0] _U435_out;
wire [15:0] _U436_in;
wire _U436_clk;
wire [15:0] _U436_out;
wire [15:0] _U437_in;
wire _U437_clk;
wire [15:0] _U437_out;
wire [15:0] _U438_in;
wire _U438_clk;
wire [15:0] _U438_out;
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
assign _U435_in = in[0];
assign _U435_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U435 (
    .in(_U435_in),
    .clk(_U435_clk),
    .out(_U435_out)
);
assign _U436_in = in[1];
assign _U436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U436 (
    .in(_U436_in),
    .clk(_U436_clk),
    .out(_U436_out)
);
assign _U437_in = in[2];
assign _U437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U437 (
    .in(_U437_in),
    .clk(_U437_clk),
    .out(_U437_out)
);
assign _U438_in = in[3];
assign _U438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(_U438_in),
    .clk(_U438_clk),
    .out(_U438_out)
);
assign _U439_in = in[4];
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign out[4] = _U439_out;
assign out[3] = _U438_out;
assign out[2] = _U437_out;
assign out[1] = _U436_out;
assign out[0] = _U435_out;
endmodule

module array_delay_U427 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U428_in;
wire _U428_clk;
wire [15:0] _U428_out;
wire [15:0] _U429_in;
wire _U429_clk;
wire [15:0] _U429_out;
wire [15:0] _U430_in;
wire _U430_clk;
wire [15:0] _U430_out;
wire [15:0] _U431_in;
wire _U431_clk;
wire [15:0] _U431_out;
wire [15:0] _U432_in;
wire _U432_clk;
wire [15:0] _U432_out;
assign _U428_in = in[0];
assign _U428_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U428_in),
    .clk(_U428_clk),
    .out(_U428_out)
);
assign _U429_in = in[1];
assign _U429_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U429 (
    .in(_U429_in),
    .clk(_U429_clk),
    .out(_U429_out)
);
assign _U430_in = in[2];
assign _U430_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U430 (
    .in(_U430_in),
    .clk(_U430_clk),
    .out(_U430_out)
);
assign _U431_in = in[3];
assign _U431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U431_in),
    .clk(_U431_clk),
    .out(_U431_out)
);
assign _U432_in = in[4];
assign _U432_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U432 (
    .in(_U432_in),
    .clk(_U432_clk),
    .out(_U432_out)
);
assign out[4] = _U432_out;
assign out[3] = _U431_out;
assign out[2] = _U430_out;
assign out[1] = _U429_out;
assign out[0] = _U428_out;
endmodule

module array_delay_U420 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire _U422_clk;
wire [15:0] _U422_out;
wire [15:0] _U423_in;
wire _U423_clk;
wire [15:0] _U423_out;
wire [15:0] _U424_in;
wire _U424_clk;
wire [15:0] _U424_out;
wire [15:0] _U425_in;
wire _U425_clk;
wire [15:0] _U425_out;
assign _U421_in = in[0];
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = in[1];
assign _U422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U422 (
    .in(_U422_in),
    .clk(_U422_clk),
    .out(_U422_out)
);
assign _U423_in = in[2];
assign _U423_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U423 (
    .in(_U423_in),
    .clk(_U423_clk),
    .out(_U423_out)
);
assign _U424_in = in[3];
assign _U424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U424 (
    .in(_U424_in),
    .clk(_U424_clk),
    .out(_U424_out)
);
assign _U425_in = in[4];
assign _U425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U425 (
    .in(_U425_in),
    .clk(_U425_clk),
    .out(_U425_out)
);
assign out[4] = _U425_out;
assign out[3] = _U424_out;
assign out[2] = _U423_out;
assign out[1] = _U422_out;
assign out[0] = _U421_out;
endmodule

module array_delay_U394 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U395_in;
wire _U395_clk;
wire [15:0] _U395_out;
wire [15:0] _U396_in;
wire _U396_clk;
wire [15:0] _U396_out;
wire [15:0] _U397_in;
wire _U397_clk;
wire [15:0] _U397_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
assign _U395_in = in[0];
assign _U395_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U395 (
    .in(_U395_in),
    .clk(_U395_clk),
    .out(_U395_out)
);
assign _U396_in = in[1];
assign _U396_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U396 (
    .in(_U396_in),
    .clk(_U396_clk),
    .out(_U396_out)
);
assign _U397_in = in[2];
assign _U397_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U397 (
    .in(_U397_in),
    .clk(_U397_clk),
    .out(_U397_out)
);
assign _U398_in = in[3];
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = in[4];
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign out[4] = _U399_out;
assign out[3] = _U398_out;
assign out[2] = _U397_out;
assign out[1] = _U396_out;
assign out[0] = _U395_out;
endmodule

module array_delay_U387 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U388_in;
wire _U388_clk;
wire [15:0] _U388_out;
wire [15:0] _U389_in;
wire _U389_clk;
wire [15:0] _U389_out;
wire [15:0] _U390_in;
wire _U390_clk;
wire [15:0] _U390_out;
wire [15:0] _U391_in;
wire _U391_clk;
wire [15:0] _U391_out;
wire [15:0] _U392_in;
wire _U392_clk;
wire [15:0] _U392_out;
assign _U388_in = in[0];
assign _U388_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U388 (
    .in(_U388_in),
    .clk(_U388_clk),
    .out(_U388_out)
);
assign _U389_in = in[1];
assign _U389_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U389 (
    .in(_U389_in),
    .clk(_U389_clk),
    .out(_U389_out)
);
assign _U390_in = in[2];
assign _U390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(_U390_in),
    .clk(_U390_clk),
    .out(_U390_out)
);
assign _U391_in = in[3];
assign _U391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U391_in),
    .clk(_U391_clk),
    .out(_U391_out)
);
assign _U392_in = in[4];
assign _U392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U392_in),
    .clk(_U392_clk),
    .out(_U392_out)
);
assign out[4] = _U392_out;
assign out[3] = _U391_out;
assign out[2] = _U390_out;
assign out[1] = _U389_out;
assign out[0] = _U388_out;
endmodule

module array_delay_U308 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire _U310_clk;
wire [15:0] _U310_out;
wire [15:0] _U311_in;
wire _U311_clk;
wire [15:0] _U311_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
wire [15:0] _U313_in;
wire _U313_clk;
wire [15:0] _U313_out;
assign _U309_in = in[0];
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = in[1];
assign _U310_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U310 (
    .in(_U310_in),
    .clk(_U310_clk),
    .out(_U310_out)
);
assign _U311_in = in[2];
assign _U311_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U311 (
    .in(_U311_in),
    .clk(_U311_clk),
    .out(_U311_out)
);
assign _U312_in = in[3];
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign _U313_in = in[4];
assign _U313_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U313 (
    .in(_U313_in),
    .clk(_U313_clk),
    .out(_U313_out)
);
assign out[4] = _U313_out;
assign out[3] = _U312_out;
assign out[2] = _U311_out;
assign out[1] = _U310_out;
assign out[0] = _U309_out;
endmodule

module array_delay_U301 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire _U303_clk;
wire [15:0] _U303_out;
wire [15:0] _U304_in;
wire _U304_clk;
wire [15:0] _U304_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
wire [15:0] _U306_in;
wire _U306_clk;
wire [15:0] _U306_out;
assign _U302_in = in[0];
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = in[1];
assign _U303_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U303 (
    .in(_U303_in),
    .clk(_U303_clk),
    .out(_U303_out)
);
assign _U304_in = in[2];
assign _U304_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U304 (
    .in(_U304_in),
    .clk(_U304_clk),
    .out(_U304_out)
);
assign _U305_in = in[3];
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign _U306_in = in[4];
assign _U306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U306_in),
    .clk(_U306_clk),
    .out(_U306_out)
);
assign out[4] = _U306_out;
assign out[3] = _U305_out;
assign out[2] = _U304_out;
assign out[1] = _U303_out;
assign out[0] = _U302_out;
endmodule

module array_delay_U294 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U295_in;
wire _U295_clk;
wire [15:0] _U295_out;
wire [15:0] _U296_in;
wire _U296_clk;
wire [15:0] _U296_out;
wire [15:0] _U297_in;
wire _U297_clk;
wire [15:0] _U297_out;
wire [15:0] _U298_in;
wire _U298_clk;
wire [15:0] _U298_out;
wire [15:0] _U299_in;
wire _U299_clk;
wire [15:0] _U299_out;
assign _U295_in = in[0];
assign _U295_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U295 (
    .in(_U295_in),
    .clk(_U295_clk),
    .out(_U295_out)
);
assign _U296_in = in[1];
assign _U296_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U296 (
    .in(_U296_in),
    .clk(_U296_clk),
    .out(_U296_out)
);
assign _U297_in = in[2];
assign _U297_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U297 (
    .in(_U297_in),
    .clk(_U297_clk),
    .out(_U297_out)
);
assign _U298_in = in[3];
assign _U298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U298 (
    .in(_U298_in),
    .clk(_U298_clk),
    .out(_U298_out)
);
assign _U299_in = in[4];
assign _U299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U299_in),
    .clk(_U299_clk),
    .out(_U299_out)
);
assign out[4] = _U299_out;
assign out[3] = _U298_out;
assign out[2] = _U297_out;
assign out[1] = _U296_out;
assign out[0] = _U295_out;
endmodule

module array_delay_U287 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U288_in;
wire _U288_clk;
wire [15:0] _U288_out;
wire [15:0] _U289_in;
wire _U289_clk;
wire [15:0] _U289_out;
wire [15:0] _U290_in;
wire _U290_clk;
wire [15:0] _U290_out;
wire [15:0] _U291_in;
wire _U291_clk;
wire [15:0] _U291_out;
wire [15:0] _U292_in;
wire _U292_clk;
wire [15:0] _U292_out;
assign _U288_in = in[0];
assign _U288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U288_in),
    .clk(_U288_clk),
    .out(_U288_out)
);
assign _U289_in = in[1];
assign _U289_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U289_in),
    .clk(_U289_clk),
    .out(_U289_out)
);
assign _U290_in = in[2];
assign _U290_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U290 (
    .in(_U290_in),
    .clk(_U290_clk),
    .out(_U290_out)
);
assign _U291_in = in[3];
assign _U291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U291 (
    .in(_U291_in),
    .clk(_U291_clk),
    .out(_U291_out)
);
assign _U292_in = in[4];
assign _U292_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U292 (
    .in(_U292_in),
    .clk(_U292_clk),
    .out(_U292_out)
);
assign out[4] = _U292_out;
assign out[3] = _U291_out;
assign out[2] = _U290_out;
assign out[1] = _U289_out;
assign out[0] = _U288_out;
endmodule

module array_delay_U280 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U281_in;
wire _U281_clk;
wire [15:0] _U281_out;
wire [15:0] _U282_in;
wire _U282_clk;
wire [15:0] _U282_out;
wire [15:0] _U283_in;
wire _U283_clk;
wire [15:0] _U283_out;
wire [15:0] _U284_in;
wire _U284_clk;
wire [15:0] _U284_out;
wire [15:0] _U285_in;
wire _U285_clk;
wire [15:0] _U285_out;
assign _U281_in = in[0];
assign _U281_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U281 (
    .in(_U281_in),
    .clk(_U281_clk),
    .out(_U281_out)
);
assign _U282_in = in[1];
assign _U282_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U282 (
    .in(_U282_in),
    .clk(_U282_clk),
    .out(_U282_out)
);
assign _U283_in = in[2];
assign _U283_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U283 (
    .in(_U283_in),
    .clk(_U283_clk),
    .out(_U283_out)
);
assign _U284_in = in[3];
assign _U284_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U284 (
    .in(_U284_in),
    .clk(_U284_clk),
    .out(_U284_out)
);
assign _U285_in = in[4];
assign _U285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(_U285_in),
    .clk(_U285_clk),
    .out(_U285_out)
);
assign out[4] = _U285_out;
assign out[3] = _U284_out;
assign out[2] = _U283_out;
assign out[1] = _U282_out;
assign out[0] = _U281_out;
endmodule

module array_delay_U273 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U274_in;
wire _U274_clk;
wire [15:0] _U274_out;
wire [15:0] _U275_in;
wire _U275_clk;
wire [15:0] _U275_out;
wire [15:0] _U276_in;
wire _U276_clk;
wire [15:0] _U276_out;
wire [15:0] _U277_in;
wire _U277_clk;
wire [15:0] _U277_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
assign _U274_in = in[0];
assign _U274_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U274 (
    .in(_U274_in),
    .clk(_U274_clk),
    .out(_U274_out)
);
assign _U275_in = in[1];
assign _U275_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U275 (
    .in(_U275_in),
    .clk(_U275_clk),
    .out(_U275_out)
);
assign _U276_in = in[2];
assign _U276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U276 (
    .in(_U276_in),
    .clk(_U276_clk),
    .out(_U276_out)
);
assign _U277_in = in[3];
assign _U277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U277 (
    .in(_U277_in),
    .clk(_U277_clk),
    .out(_U277_out)
);
assign _U278_in = in[4];
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign out[4] = _U278_out;
assign out[3] = _U277_out;
assign out[2] = _U276_out;
assign out[1] = _U275_out;
assign out[0] = _U274_out;
endmodule

module array_delay_U266 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire _U268_clk;
wire [15:0] _U268_out;
wire [15:0] _U269_in;
wire _U269_clk;
wire [15:0] _U269_out;
wire [15:0] _U270_in;
wire _U270_clk;
wire [15:0] _U270_out;
wire [15:0] _U271_in;
wire _U271_clk;
wire [15:0] _U271_out;
assign _U267_in = in[0];
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = in[1];
assign _U268_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U268 (
    .in(_U268_in),
    .clk(_U268_clk),
    .out(_U268_out)
);
assign _U269_in = in[2];
assign _U269_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U269 (
    .in(_U269_in),
    .clk(_U269_clk),
    .out(_U269_out)
);
assign _U270_in = in[3];
assign _U270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(_U270_in),
    .clk(_U270_clk),
    .out(_U270_out)
);
assign _U271_in = in[4];
assign _U271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U271_in),
    .clk(_U271_clk),
    .out(_U271_out)
);
assign out[4] = _U271_out;
assign out[3] = _U270_out;
assign out[2] = _U269_out;
assign out[1] = _U268_out;
assign out[0] = _U267_out;
endmodule

module array_delay_U259 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U260_in;
wire _U260_clk;
wire [15:0] _U260_out;
wire [15:0] _U261_in;
wire _U261_clk;
wire [15:0] _U261_out;
wire [15:0] _U262_in;
wire _U262_clk;
wire [15:0] _U262_out;
wire [15:0] _U263_in;
wire _U263_clk;
wire [15:0] _U263_out;
wire [15:0] _U264_in;
wire _U264_clk;
wire [15:0] _U264_out;
assign _U260_in = in[0];
assign _U260_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U260_in),
    .clk(_U260_clk),
    .out(_U260_out)
);
assign _U261_in = in[1];
assign _U261_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U261 (
    .in(_U261_in),
    .clk(_U261_clk),
    .out(_U261_out)
);
assign _U262_in = in[2];
assign _U262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U262 (
    .in(_U262_in),
    .clk(_U262_clk),
    .out(_U262_out)
);
assign _U263_in = in[3];
assign _U263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U263 (
    .in(_U263_in),
    .clk(_U263_clk),
    .out(_U263_out)
);
assign _U264_in = in[4];
assign _U264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U264_in),
    .clk(_U264_clk),
    .out(_U264_out)
);
assign out[4] = _U264_out;
assign out[3] = _U263_out;
assign out[2] = _U262_out;
assign out[1] = _U261_out;
assign out[0] = _U260_out;
endmodule

module array_delay_U252 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U253_in;
wire _U253_clk;
wire [15:0] _U253_out;
wire [15:0] _U254_in;
wire _U254_clk;
wire [15:0] _U254_out;
wire [15:0] _U255_in;
wire _U255_clk;
wire [15:0] _U255_out;
wire [15:0] _U256_in;
wire _U256_clk;
wire [15:0] _U256_out;
wire [15:0] _U257_in;
wire _U257_clk;
wire [15:0] _U257_out;
assign _U253_in = in[0];
assign _U253_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U253 (
    .in(_U253_in),
    .clk(_U253_clk),
    .out(_U253_out)
);
assign _U254_in = in[1];
assign _U254_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U254 (
    .in(_U254_in),
    .clk(_U254_clk),
    .out(_U254_out)
);
assign _U255_in = in[2];
assign _U255_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U255 (
    .in(_U255_in),
    .clk(_U255_clk),
    .out(_U255_out)
);
assign _U256_in = in[3];
assign _U256_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U256 (
    .in(_U256_in),
    .clk(_U256_clk),
    .out(_U256_out)
);
assign _U257_in = in[4];
assign _U257_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U257 (
    .in(_U257_in),
    .clk(_U257_clk),
    .out(_U257_out)
);
assign out[4] = _U257_out;
assign out[3] = _U256_out;
assign out[2] = _U255_out;
assign out[1] = _U254_out;
assign out[0] = _U253_out;
endmodule

module array_delay_U245 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U246_in;
wire _U246_clk;
wire [15:0] _U246_out;
wire [15:0] _U247_in;
wire _U247_clk;
wire [15:0] _U247_out;
wire [15:0] _U248_in;
wire _U248_clk;
wire [15:0] _U248_out;
wire [15:0] _U249_in;
wire _U249_clk;
wire [15:0] _U249_out;
wire [15:0] _U250_in;
wire _U250_clk;
wire [15:0] _U250_out;
assign _U246_in = in[0];
assign _U246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(_U246_in),
    .clk(_U246_clk),
    .out(_U246_out)
);
assign _U247_in = in[1];
assign _U247_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U247 (
    .in(_U247_in),
    .clk(_U247_clk),
    .out(_U247_out)
);
assign _U248_in = in[2];
assign _U248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U248 (
    .in(_U248_in),
    .clk(_U248_clk),
    .out(_U248_out)
);
assign _U249_in = in[3];
assign _U249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U249 (
    .in(_U249_in),
    .clk(_U249_clk),
    .out(_U249_out)
);
assign _U250_in = in[4];
assign _U250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U250 (
    .in(_U250_in),
    .clk(_U250_clk),
    .out(_U250_out)
);
assign out[4] = _U250_out;
assign out[3] = _U249_out;
assign out[2] = _U248_out;
assign out[1] = _U247_out;
assign out[0] = _U246_out;
endmodule

module array_delay_U238 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U239_in;
wire _U239_clk;
wire [15:0] _U239_out;
wire [15:0] _U240_in;
wire _U240_clk;
wire [15:0] _U240_out;
wire [15:0] _U241_in;
wire _U241_clk;
wire [15:0] _U241_out;
wire [15:0] _U242_in;
wire _U242_clk;
wire [15:0] _U242_out;
wire [15:0] _U243_in;
wire _U243_clk;
wire [15:0] _U243_out;
assign _U239_in = in[0];
assign _U239_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U239 (
    .in(_U239_in),
    .clk(_U239_clk),
    .out(_U239_out)
);
assign _U240_in = in[1];
assign _U240_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U240 (
    .in(_U240_in),
    .clk(_U240_clk),
    .out(_U240_out)
);
assign _U241_in = in[2];
assign _U241_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U241 (
    .in(_U241_in),
    .clk(_U241_clk),
    .out(_U241_out)
);
assign _U242_in = in[3];
assign _U242_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U242 (
    .in(_U242_in),
    .clk(_U242_clk),
    .out(_U242_out)
);
assign _U243_in = in[4];
assign _U243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U243_in),
    .clk(_U243_clk),
    .out(_U243_out)
);
assign out[4] = _U243_out;
assign out[3] = _U242_out;
assign out[2] = _U241_out;
assign out[1] = _U240_out;
assign out[0] = _U239_out;
endmodule

module array_delay_U231 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
wire [15:0] _U233_in;
wire _U233_clk;
wire [15:0] _U233_out;
wire [15:0] _U234_in;
wire _U234_clk;
wire [15:0] _U234_out;
wire [15:0] _U235_in;
wire _U235_clk;
wire [15:0] _U235_out;
wire [15:0] _U236_in;
wire _U236_clk;
wire [15:0] _U236_out;
assign _U232_in = in[0];
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign _U233_in = in[1];
assign _U233_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U233 (
    .in(_U233_in),
    .clk(_U233_clk),
    .out(_U233_out)
);
assign _U234_in = in[2];
assign _U234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U234 (
    .in(_U234_in),
    .clk(_U234_clk),
    .out(_U234_out)
);
assign _U235_in = in[3];
assign _U235_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U235 (
    .in(_U235_in),
    .clk(_U235_clk),
    .out(_U235_out)
);
assign _U236_in = in[4];
assign _U236_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U236 (
    .in(_U236_in),
    .clk(_U236_clk),
    .out(_U236_out)
);
assign out[4] = _U236_out;
assign out[3] = _U235_out;
assign out[2] = _U234_out;
assign out[1] = _U233_out;
assign out[0] = _U232_out;
endmodule

module array_delay_U224 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire _U228_clk;
wire [15:0] _U228_out;
wire [15:0] _U229_in;
wire _U229_clk;
wire [15:0] _U229_out;
assign _U225_in = in[0];
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = in[1];
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = in[2];
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = in[3];
assign _U228_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U228 (
    .in(_U228_in),
    .clk(_U228_clk),
    .out(_U228_out)
);
assign _U229_in = in[4];
assign _U229_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U229 (
    .in(_U229_in),
    .clk(_U229_clk),
    .out(_U229_out)
);
assign out[4] = _U229_out;
assign out[3] = _U228_out;
assign out[2] = _U227_out;
assign out[1] = _U226_out;
assign out[0] = _U225_out;
endmodule

module array_delay_U217 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
wire [15:0] _U219_in;
wire _U219_clk;
wire [15:0] _U219_out;
wire [15:0] _U220_in;
wire _U220_clk;
wire [15:0] _U220_out;
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
assign _U218_in = in[0];
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign _U219_in = in[1];
assign _U219_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U219_in),
    .clk(_U219_clk),
    .out(_U219_out)
);
assign _U220_in = in[2];
assign _U220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U220_in),
    .clk(_U220_clk),
    .out(_U220_out)
);
assign _U221_in = in[3];
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign _U222_in = in[4];
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign out[4] = _U222_out;
assign out[3] = _U221_out;
assign out[2] = _U220_out;
assign out[1] = _U219_out;
assign out[0] = _U218_out;
endmodule

module array_delay_U210 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U211_in;
wire _U211_clk;
wire [15:0] _U211_out;
wire [15:0] _U212_in;
wire _U212_clk;
wire [15:0] _U212_out;
wire [15:0] _U213_in;
wire _U213_clk;
wire [15:0] _U213_out;
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire _U215_clk;
wire [15:0] _U215_out;
assign _U211_in = in[0];
assign _U211_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U211 (
    .in(_U211_in),
    .clk(_U211_clk),
    .out(_U211_out)
);
assign _U212_in = in[1];
assign _U212_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U212 (
    .in(_U212_in),
    .clk(_U212_clk),
    .out(_U212_out)
);
assign _U213_in = in[2];
assign _U213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(_U213_in),
    .clk(_U213_clk),
    .out(_U213_out)
);
assign _U214_in = in[3];
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = in[4];
assign _U215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(_U215_in),
    .clk(_U215_clk),
    .out(_U215_out)
);
assign out[4] = _U215_out;
assign out[3] = _U214_out;
assign out[2] = _U213_out;
assign out[1] = _U212_out;
assign out[0] = _U211_out;
endmodule

module array_delay_U203 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U205_in;
wire _U205_clk;
wire [15:0] _U205_out;
wire [15:0] _U206_in;
wire _U206_clk;
wire [15:0] _U206_out;
wire [15:0] _U207_in;
wire _U207_clk;
wire [15:0] _U207_out;
wire [15:0] _U208_in;
wire _U208_clk;
wire [15:0] _U208_out;
assign _U204_in = in[0];
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U205_in = in[1];
assign _U205_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U205 (
    .in(_U205_in),
    .clk(_U205_clk),
    .out(_U205_out)
);
assign _U206_in = in[2];
assign _U206_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U206 (
    .in(_U206_in),
    .clk(_U206_clk),
    .out(_U206_out)
);
assign _U207_in = in[3];
assign _U207_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U207 (
    .in(_U207_in),
    .clk(_U207_clk),
    .out(_U207_out)
);
assign _U208_in = in[4];
assign _U208_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U208 (
    .in(_U208_in),
    .clk(_U208_clk),
    .out(_U208_out)
);
assign out[4] = _U208_out;
assign out[3] = _U207_out;
assign out[2] = _U206_out;
assign out[1] = _U205_out;
assign out[0] = _U204_out;
endmodule

module array_delay_U196 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U197_in;
wire _U197_clk;
wire [15:0] _U197_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire _U199_clk;
wire [15:0] _U199_out;
wire [15:0] _U200_in;
wire _U200_clk;
wire [15:0] _U200_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
assign _U197_in = in[0];
assign _U197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U197 (
    .in(_U197_in),
    .clk(_U197_clk),
    .out(_U197_out)
);
assign _U198_in = in[1];
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = in[2];
assign _U199_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U199 (
    .in(_U199_in),
    .clk(_U199_clk),
    .out(_U199_out)
);
assign _U200_in = in[3];
assign _U200_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U200 (
    .in(_U200_in),
    .clk(_U200_clk),
    .out(_U200_out)
);
assign _U201_in = in[4];
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign out[4] = _U201_out;
assign out[3] = _U200_out;
assign out[2] = _U199_out;
assign out[1] = _U198_out;
assign out[0] = _U197_out;
endmodule

module array_delay_U170 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire _U172_clk;
wire [15:0] _U172_out;
wire [15:0] _U173_in;
wire _U173_clk;
wire [15:0] _U173_out;
wire [15:0] _U174_in;
wire _U174_clk;
wire [15:0] _U174_out;
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
assign _U171_in = in[0];
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = in[1];
assign _U172_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U172 (
    .in(_U172_in),
    .clk(_U172_clk),
    .out(_U172_out)
);
assign _U173_in = in[2];
assign _U173_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U173 (
    .in(_U173_in),
    .clk(_U173_clk),
    .out(_U173_out)
);
assign _U174_in = in[3];
assign _U174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(_U174_in),
    .clk(_U174_clk),
    .out(_U174_out)
);
assign _U175_in = in[4];
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign out[4] = _U175_out;
assign out[3] = _U174_out;
assign out[2] = _U173_out;
assign out[1] = _U172_out;
assign out[0] = _U171_out;
endmodule

module array_delay_U163 (
    input clk,
    input [15:0] in [4:0],
    output [15:0] out [4:0]
);
wire [15:0] _U164_in;
wire _U164_clk;
wire [15:0] _U164_out;
wire [15:0] _U165_in;
wire _U165_clk;
wire [15:0] _U165_out;
wire [15:0] _U166_in;
wire _U166_clk;
wire [15:0] _U166_out;
wire [15:0] _U167_in;
wire _U167_clk;
wire [15:0] _U167_out;
wire [15:0] _U168_in;
wire _U168_clk;
wire [15:0] _U168_out;
assign _U164_in = in[0];
assign _U164_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U164 (
    .in(_U164_in),
    .clk(_U164_clk),
    .out(_U164_out)
);
assign _U165_in = in[1];
assign _U165_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U165 (
    .in(_U165_in),
    .clk(_U165_clk),
    .out(_U165_out)
);
assign _U166_in = in[2];
assign _U166_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(_U166_in),
    .clk(_U166_clk),
    .out(_U166_out)
);
assign _U167_in = in[3];
assign _U167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U167_in),
    .clk(_U167_clk),
    .out(_U167_out)
);
assign _U168_in = in[4];
assign _U168_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U168 (
    .in(_U168_in),
    .clk(_U168_clk),
    .out(_U168_out)
);
assign out[4] = _U168_out;
assign out[3] = _U167_out;
assign out[2] = _U166_out;
assign out[1] = _U165_out;
assign out[0] = _U164_out;
endmodule

module array_delay_U121 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U122_in;
wire _U122_clk;
wire [15:0] _U122_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire _U124_clk;
wire [15:0] _U124_out;
wire [15:0] _U125_in;
wire _U125_clk;
wire [15:0] _U125_out;
assign _U122_in = in[0];
assign _U122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U122 (
    .in(_U122_in),
    .clk(_U122_clk),
    .out(_U122_out)
);
assign _U123_in = in[1];
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = in[2];
assign _U124_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U124 (
    .in(_U124_in),
    .clk(_U124_clk),
    .out(_U124_out)
);
assign _U125_in = in[3];
assign _U125_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U125 (
    .in(_U125_in),
    .clk(_U125_clk),
    .out(_U125_out)
);
assign out[3] = _U125_out;
assign out[2] = _U124_out;
assign out[1] = _U123_out;
assign out[0] = _U122_out;
endmodule

module array_delay_U115 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U116_in;
wire _U116_clk;
wire [15:0] _U116_out;
wire [15:0] _U117_in;
wire _U117_clk;
wire [15:0] _U117_out;
wire [15:0] _U118_in;
wire _U118_clk;
wire [15:0] _U118_out;
wire [15:0] _U119_in;
wire _U119_clk;
wire [15:0] _U119_out;
assign _U116_in = in[0];
assign _U116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U116_in),
    .clk(_U116_clk),
    .out(_U116_out)
);
assign _U117_in = in[1];
assign _U117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U117 (
    .in(_U117_in),
    .clk(_U117_clk),
    .out(_U117_out)
);
assign _U118_in = in[2];
assign _U118_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U118 (
    .in(_U118_in),
    .clk(_U118_clk),
    .out(_U118_out)
);
assign _U119_in = in[3];
assign _U119_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U119 (
    .in(_U119_in),
    .clk(_U119_clk),
    .out(_U119_out)
);
assign out[3] = _U119_out;
assign out[2] = _U118_out;
assign out[1] = _U117_out;
assign out[0] = _U116_out;
endmodule

module array_delay_U105 (
    input clk,
    input [15:0] in [3:0],
    output [15:0] out [3:0]
);
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire _U108_clk;
wire [15:0] _U108_out;
wire [15:0] _U109_in;
wire _U109_clk;
wire [15:0] _U109_out;
assign _U106_in = in[0];
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = in[1];
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = in[2];
assign _U108_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U108 (
    .in(_U108_in),
    .clk(_U108_clk),
    .out(_U108_out)
);
assign _U109_in = in[3];
assign _U109_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U109 (
    .in(_U109_in),
    .clk(_U109_clk),
    .out(_U109_out)
);
assign out[3] = _U109_out;
assign out[2] = _U108_out;
assign out[1] = _U107_out;
assign out[0] = _U106_out;
endmodule

module aff__U727 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h010e * d[1])))) + (16'(16'h0009 * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h0001);
endmodule

module affine_controller__U726 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U727 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001d;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001d;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0007;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U70 (
    output [15:0] out,
    input [15:0] d [3:0]
);
assign out = 16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h032c * d[1])))) + (16'(16'h001d * d[2])))) + (16'(16'h0001 * d[3])))) + 16'h7d21);
endmodule

module affine_controller__U69 (
    input clk,
    output valid,
    output [15:0] d [3:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [3:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U70 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = ((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = (1'b1 & d_2_at_max_out) & d_3_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 & d_3_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign valid = cmp_time_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U539 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U538 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U539 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U47 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U46 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U47 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U351 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U350 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U351 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U315 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0051 * d[1])))) + (16'(16'h001b * d[2])))) + (16'(16'h0009 * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h0002);
endmodule

module affine_controller__U314 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U315 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h0002;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h0007;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U24 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U23 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U24 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U127 (
    output [15:0] out,
    input [15:0] d [4:0]
);
assign out = 16'((16'((16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h0f18 * d[1])))) + (16'(16'h0508 * d[2])))) + (16'(16'h002e * d[3])))) + (16'(16'h0001 * d[4])))) + 16'h1f49);
endmodule

module affine_controller__U126 (
    input clk,
    output valid,
    output [15:0] d [4:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [4:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
wire d_3_at_max_out;
wire [15:0] d_3_reg_in;
wire d_3_reg_clk;
wire [15:0] d_3_reg_out;
wire d_3_reg_en;
wire d_4_at_max_out;
wire [15:0] d_4_reg_in;
wire d_4_reg_clk;
wire [15:0] d_4_reg_out;
wire d_4_reg_en;
assign affine_func_d[4] = d_4_reg_out;
assign affine_func_d[3] = d_3_reg_out;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U127 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (((1'b1 & d_1_at_max_out) & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h0002;
assign d_1_reg_in = ((1'b1 & d_2_at_max_out) & d_3_at_max_out) & d_4_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h0002;
assign d_2_reg_in = (1'b1 & d_3_at_max_out) & d_4_at_max_out ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign d_3_at_max_out = d_3_reg_out == 16'h001b;
assign d_3_reg_in = 1'b1 & d_4_at_max_out ? d_3_at_max_out ? 16'h0000 : 16'(d_3_reg_out + 16'h0001) : d_3_reg_out;
assign d_3_reg_clk = clk;
assign d_3_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_3_reg (
    .in(d_3_reg_in),
    .clk(d_3_reg_clk),
    .out(d_3_reg_out),
    .en(d_3_reg_en)
);
assign d_4_at_max_out = d_4_reg_out == 16'h001b;
assign d_4_reg_in = 1'b1 ? d_4_at_max_out ? 16'h0000 : 16'(d_4_reg_out + 16'h0001) : d_4_reg_out;
assign d_4_reg_clk = clk;
assign d_4_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_4_reg (
    .in(d_4_reg_in),
    .clk(d_4_reg_clk),
    .out(d_4_reg_out),
    .en(d_4_reg_en)
);
assign valid = cmp_time_out;
assign d[4] = d_4_reg_out;
assign d[3] = d_3_reg_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module aff__U1 (
    output [15:0] out,
    input [15:0] d [2:0]
);
assign out = 16'((16'((16'((16'(16'h0000 * d[0])) + (16'(16'h001d * d[1])))) + (16'(16'h0001 * d[2])))) + 16'h0002);
endmodule

module affine_controller__U0 (
    input clk,
    output valid,
    output [15:0] d [2:0]
);
wire [15:0] affine_func_out;
wire [15:0] affine_func_d [2:0];
wire cmp_time_out;
wire [15:0] cycle_time_in;
wire cycle_time_clk;
wire [15:0] cycle_time_out;
wire [15:0] d_0_reg_in;
wire d_0_reg_clk;
wire [15:0] d_0_reg_out;
wire d_0_reg_en;
wire d_1_at_max_out;
wire [15:0] d_1_reg_in;
wire d_1_reg_clk;
wire [15:0] d_1_reg_out;
wire d_1_reg_en;
wire d_2_at_max_out;
wire [15:0] d_2_reg_in;
wire d_2_reg_clk;
wire [15:0] d_2_reg_out;
wire d_2_reg_en;
assign affine_func_d[2] = d_2_reg_out;
assign affine_func_d[1] = d_1_reg_out;
assign affine_func_d[0] = d_0_reg_out;
aff__U1 affine_func (
    .out(affine_func_out),
    .d(affine_func_d)
);
assign cmp_time_out = (16'(affine_func_out - cycle_time_out)) == 16'h0000;
assign cycle_time_in = 16'(cycle_time_out + 16'h0001);
assign cycle_time_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) cycle_time (
    .in(cycle_time_in),
    .clk(cycle_time_clk),
    .out(cycle_time_out)
);
assign d_0_reg_in = (1'b1 & d_1_at_max_out) & d_2_at_max_out ? d_0_reg_out == 16'h0000 ? 16'h0000 : 16'(d_0_reg_out + 16'h0001) : d_0_reg_out;
assign d_0_reg_clk = clk;
assign d_0_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_0_reg (
    .in(d_0_reg_in),
    .clk(d_0_reg_clk),
    .out(d_0_reg_out),
    .en(d_0_reg_en)
);
assign d_1_at_max_out = d_1_reg_out == 16'h001b;
assign d_1_reg_in = 1'b1 & d_2_at_max_out ? d_1_at_max_out ? 16'h0000 : 16'(d_1_reg_out + 16'h0001) : d_1_reg_out;
assign d_1_reg_clk = clk;
assign d_1_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_1_reg (
    .in(d_1_reg_in),
    .clk(d_1_reg_clk),
    .out(d_1_reg_out),
    .en(d_1_reg_en)
);
assign d_2_at_max_out = d_2_reg_out == 16'h001b;
assign d_2_reg_in = 1'b1 ? d_2_at_max_out ? 16'h0000 : 16'(d_2_reg_out + 16'h0001) : d_2_reg_out;
assign d_2_reg_clk = clk;
assign d_2_reg_en = cmp_time_out;
mantle_reg__has_clrFalse__has_enTrue__has_rstFalse__width16 #(
    .init(16'h0000)
) d_2_reg (
    .in(d_2_reg_in),
    .clk(d_2_reg_clk),
    .out(d_2_reg_out),
    .en(d_2_reg_en)
);
assign valid = cmp_time_out;
assign d[2] = d_2_reg_out;
assign d[1] = d_1_reg_out;
assign d[0] = d_0_reg_out;
endmodule

module _U97_pt__U98 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U8_pt__U9 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U86_pt__U87 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U76_pt__U77 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U73_pt__U74 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U71_pt__U72 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U6_pt__U7 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_output_stencil_pipelined (
    output [15:0] out_hw_output_stencil,
    input [15:0] in0_conv_stencil [0:0]
);
wire [15:0] _U6_in;
assign _U6_in = in0_conv_stencil[0];
_U6_pt__U7 _U6 (
    .in(_U6_in),
    .out(out_hw_output_stencil)
);
endmodule

module cu_op_hcompute_hw_output_stencil (
    input clk,
    input [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0],
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_output_stencil;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
hcompute_hw_output_stencil_pipelined inner_compute (
    .out_hw_output_stencil(inner_compute_out_hw_output_stencil),
    .in0_conv_stencil(inner_compute_in0_conv_stencil)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = inner_compute_out_hw_output_stencil;
endmodule

module _U69_pt__U70 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U67_pt__U68 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U64_pt__U65 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U613_pt__U614 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_input_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_input_global_wrapper_stencil,
    input [15:0] in0_hw_input_stencil [0:0]
);
wire [15:0] _U613_in;
assign _U613_in = in0_hw_input_stencil[0];
_U613_pt__U614 _U613 (
    .in(_U613_in),
    .out(out_hw_input_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_input_global_wrapper_stencil (
    input clk,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_input_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_input_stencil [0:0];
assign inner_compute_in0_hw_input_stencil[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
hcompute_hw_input_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_input_global_wrapper_stencil(inner_compute_out_hw_input_global_wrapper_stencil),
    .in0_hw_input_stencil(inner_compute_in0_hw_input_stencil)
);
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = inner_compute_out_hw_input_global_wrapper_stencil;
endmodule

module _U604_pt__U605 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U595_pt__U596 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U587_pt__U588 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U579_pt__U580 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U572_pt__U573 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U565_pt__U566 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U559_pt__U560 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U553_pt__U554 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U548_pt__U549 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U543_pt__U544 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U539_pt__U540 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U535_pt__U536 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U532_pt__U533 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U52_pt__U53 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U529_pt__U530 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U527_pt__U528 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U525_pt__U526 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U509_pt__U510 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U506_pt__U507 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U502_pt__U503 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U4_pt__U5 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_2_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U4_in;
assign _U4_in = 16'h0000;
_U4_pt__U5 _U4 (
    .in(_U4_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_2 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_2_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U499_pt__U500 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U493_pt__U494 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U490_pt__U491 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U482_pt__U483 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U47_pt__U48 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U479_pt__U480 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U469_pt__U470 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U466_pt__U467 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U454_pt__U455 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U451_pt__U452 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U44_pt__U45 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U448_pt__U449 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U434_pt__U435 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U432_pt__U433 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U429_pt__U430 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U41_pt__U42 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U412_pt__U413 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_3_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U412_in;
wire [15:0] _U412_out;
wire [15:0] _U414_in;
wire _U414_clk;
wire [15:0] _U414_out;
wire [15:0] _U415_in;
wire _U415_clk;
wire [15:0] _U415_out;
wire [15:0] _U416_in;
wire _U416_clk;
wire [15:0] _U416_out;
wire [15:0] _U417_in;
wire _U417_clk;
wire [15:0] _U417_out;
wire [15:0] _U418_in;
wire _U418_clk;
wire [15:0] _U418_out;
wire [15:0] _U419_in;
wire _U419_clk;
wire [15:0] _U419_out;
wire [15:0] _U420_in;
wire _U420_clk;
wire [15:0] _U420_out;
wire [15:0] _U421_in;
wire _U421_clk;
wire [15:0] _U421_out;
wire [15:0] _U422_in;
wire _U422_clk;
wire [15:0] _U422_out;
wire [15:0] _U423_in;
wire _U423_clk;
wire [15:0] _U423_out;
wire [15:0] _U424_in;
wire _U424_clk;
wire [15:0] _U424_out;
wire [15:0] _U425_in;
wire _U425_clk;
wire [15:0] _U425_out;
wire [15:0] _U426_in;
wire _U426_clk;
wire [15:0] _U426_out;
wire [15:0] _U427_in;
wire _U427_clk;
wire [15:0] _U427_out;
wire [15:0] _U428_in;
wire _U428_clk;
wire [15:0] _U428_out;
wire [15:0] _U429_in;
wire [15:0] _U429_out;
wire [15:0] _U431_in;
wire _U431_clk;
wire [15:0] _U431_out;
wire [15:0] _U432_in;
wire [15:0] _U434_in;
wire [15:0] _U434_out;
wire [15:0] _U436_in;
wire _U436_clk;
wire [15:0] _U436_out;
wire [15:0] _U437_in;
wire _U437_clk;
wire [15:0] _U437_out;
wire [15:0] _U438_in;
wire _U438_clk;
wire [15:0] _U438_out;
wire [15:0] _U439_in;
wire _U439_clk;
wire [15:0] _U439_out;
wire [15:0] _U440_in;
wire _U440_clk;
wire [15:0] _U440_out;
wire [15:0] _U441_in;
wire _U441_clk;
wire [15:0] _U441_out;
wire [15:0] _U442_in;
wire _U442_clk;
wire [15:0] _U442_out;
wire [15:0] _U443_in;
wire _U443_clk;
wire [15:0] _U443_out;
wire [15:0] _U444_in;
wire _U444_clk;
wire [15:0] _U444_out;
wire [15:0] _U445_in;
wire _U445_clk;
wire [15:0] _U445_out;
wire [15:0] _U446_in;
wire _U446_clk;
wire [15:0] _U446_out;
wire [15:0] _U447_in;
wire _U447_clk;
wire [15:0] _U447_out;
wire [15:0] _U448_in;
wire [15:0] _U448_out;
wire [15:0] _U450_in;
wire _U450_clk;
wire [15:0] _U450_out;
wire [15:0] _U451_in;
wire [15:0] _U451_out;
wire [15:0] _U453_in;
wire _U453_clk;
wire [15:0] _U453_out;
wire [15:0] _U454_in;
wire [15:0] _U454_out;
wire [15:0] _U456_in;
wire _U456_clk;
wire [15:0] _U456_out;
wire [15:0] _U457_in;
wire _U457_clk;
wire [15:0] _U457_out;
wire [15:0] _U458_in;
wire _U458_clk;
wire [15:0] _U458_out;
wire [15:0] _U459_in;
wire _U459_clk;
wire [15:0] _U459_out;
wire [15:0] _U460_in;
wire _U460_clk;
wire [15:0] _U460_out;
wire [15:0] _U461_in;
wire _U461_clk;
wire [15:0] _U461_out;
wire [15:0] _U462_in;
wire _U462_clk;
wire [15:0] _U462_out;
wire [15:0] _U463_in;
wire _U463_clk;
wire [15:0] _U463_out;
wire [15:0] _U464_in;
wire _U464_clk;
wire [15:0] _U464_out;
wire [15:0] _U465_in;
wire _U465_clk;
wire [15:0] _U465_out;
wire [15:0] _U466_in;
wire [15:0] _U466_out;
wire [15:0] _U468_in;
wire _U468_clk;
wire [15:0] _U468_out;
wire [15:0] _U469_in;
wire [15:0] _U469_out;
wire [15:0] _U471_in;
wire _U471_clk;
wire [15:0] _U471_out;
wire [15:0] _U472_in;
wire _U472_clk;
wire [15:0] _U472_out;
wire [15:0] _U473_in;
wire _U473_clk;
wire [15:0] _U473_out;
wire [15:0] _U474_in;
wire _U474_clk;
wire [15:0] _U474_out;
wire [15:0] _U475_in;
wire _U475_clk;
wire [15:0] _U475_out;
wire [15:0] _U476_in;
wire _U476_clk;
wire [15:0] _U476_out;
wire [15:0] _U477_in;
wire _U477_clk;
wire [15:0] _U477_out;
wire [15:0] _U478_in;
wire _U478_clk;
wire [15:0] _U478_out;
wire [15:0] _U479_in;
wire [15:0] _U479_out;
wire [15:0] _U481_in;
wire _U481_clk;
wire [15:0] _U481_out;
wire [15:0] _U482_in;
wire [15:0] _U482_out;
wire [15:0] _U484_in;
wire _U484_clk;
wire [15:0] _U484_out;
wire [15:0] _U485_in;
wire _U485_clk;
wire [15:0] _U485_out;
wire [15:0] _U486_in;
wire _U486_clk;
wire [15:0] _U486_out;
wire [15:0] _U487_in;
wire _U487_clk;
wire [15:0] _U487_out;
wire [15:0] _U488_in;
wire _U488_clk;
wire [15:0] _U488_out;
wire [15:0] _U489_in;
wire _U489_clk;
wire [15:0] _U489_out;
wire [15:0] _U490_in;
wire [15:0] _U490_out;
wire [15:0] _U492_in;
wire _U492_clk;
wire [15:0] _U492_out;
wire [15:0] _U493_in;
wire [15:0] _U493_out;
wire [15:0] _U495_in;
wire _U495_clk;
wire [15:0] _U495_out;
wire [15:0] _U496_in;
wire _U496_clk;
wire [15:0] _U496_out;
wire [15:0] _U497_in;
wire _U497_clk;
wire [15:0] _U497_out;
wire [15:0] _U498_in;
wire _U498_clk;
wire [15:0] _U498_out;
wire [15:0] _U499_in;
wire [15:0] _U499_out;
wire [15:0] _U501_in;
wire _U501_clk;
wire [15:0] _U501_out;
wire [15:0] _U502_in;
wire [15:0] _U502_out;
wire [15:0] _U504_in;
wire _U504_clk;
wire [15:0] _U504_out;
wire [15:0] _U505_in;
wire _U505_clk;
wire [15:0] _U505_out;
wire [15:0] _U506_in;
wire [15:0] _U506_out;
wire [15:0] _U508_in;
wire _U508_clk;
wire [15:0] _U508_out;
wire [15:0] _U509_in;
wire [15:0] _U509_out;
wire [15:0] _U511_in;
wire _U511_clk;
wire [15:0] _U511_out;
wire [15:0] _U512_in;
wire _U512_clk;
wire [15:0] _U512_out;
wire [15:0] _U513_in;
wire _U513_clk;
wire [15:0] _U513_out;
wire [15:0] _U514_in;
wire _U514_clk;
wire [15:0] _U514_out;
wire [15:0] _U515_in;
wire _U515_clk;
wire [15:0] _U515_out;
wire [15:0] _U516_in;
wire _U516_clk;
wire [15:0] _U516_out;
wire [15:0] _U517_in;
wire _U517_clk;
wire [15:0] _U517_out;
wire [15:0] _U518_in;
wire _U518_clk;
wire [15:0] _U518_out;
wire [15:0] _U519_in;
wire _U519_clk;
wire [15:0] _U519_out;
wire [15:0] _U520_in;
wire _U520_clk;
wire [15:0] _U520_out;
wire [15:0] _U521_in;
wire _U521_clk;
wire [15:0] _U521_out;
wire [15:0] _U522_in;
wire _U522_clk;
wire [15:0] _U522_out;
wire [15:0] _U523_in;
wire _U523_clk;
wire [15:0] _U523_out;
wire [15:0] _U524_in;
wire _U524_clk;
wire [15:0] _U524_out;
wire [15:0] _U525_in;
wire [15:0] _U525_out;
wire [15:0] _U527_in;
wire [15:0] _U527_out;
wire [15:0] _U529_in;
wire [15:0] _U529_out;
wire [15:0] _U531_in;
wire _U531_clk;
wire [15:0] _U531_out;
wire [15:0] _U532_in;
wire [15:0] _U532_out;
wire [15:0] _U534_in;
wire _U534_clk;
wire [15:0] _U534_out;
wire [15:0] _U535_in;
wire [15:0] _U535_out;
wire [15:0] _U537_in;
wire _U537_clk;
wire [15:0] _U537_out;
wire [15:0] _U538_in;
wire _U538_clk;
wire [15:0] _U538_out;
wire [15:0] _U539_in;
wire [15:0] _U539_out;
wire [15:0] _U541_in;
wire _U541_clk;
wire [15:0] _U541_out;
wire [15:0] _U542_in;
wire _U542_clk;
wire [15:0] _U542_out;
wire [15:0] _U543_in;
wire [15:0] _U543_out;
wire [15:0] _U545_in;
wire _U545_clk;
wire [15:0] _U545_out;
wire [15:0] _U546_in;
wire _U546_clk;
wire [15:0] _U546_out;
wire [15:0] _U547_in;
wire _U547_clk;
wire [15:0] _U547_out;
wire [15:0] _U548_in;
wire [15:0] _U548_out;
wire [15:0] _U550_in;
wire _U550_clk;
wire [15:0] _U550_out;
wire [15:0] _U551_in;
wire _U551_clk;
wire [15:0] _U551_out;
wire [15:0] _U552_in;
wire _U552_clk;
wire [15:0] _U552_out;
wire [15:0] _U553_in;
wire [15:0] _U553_out;
wire [15:0] _U555_in;
wire _U555_clk;
wire [15:0] _U555_out;
wire [15:0] _U556_in;
wire _U556_clk;
wire [15:0] _U556_out;
wire [15:0] _U557_in;
wire _U557_clk;
wire [15:0] _U557_out;
wire [15:0] _U558_in;
wire _U558_clk;
wire [15:0] _U558_out;
wire [15:0] _U559_in;
wire [15:0] _U559_out;
wire [15:0] _U561_in;
wire _U561_clk;
wire [15:0] _U561_out;
wire [15:0] _U562_in;
wire _U562_clk;
wire [15:0] _U562_out;
wire [15:0] _U563_in;
wire _U563_clk;
wire [15:0] _U563_out;
wire [15:0] _U564_in;
wire _U564_clk;
wire [15:0] _U564_out;
wire [15:0] _U565_in;
wire [15:0] _U565_out;
wire [15:0] _U567_in;
wire _U567_clk;
wire [15:0] _U567_out;
wire [15:0] _U568_in;
wire _U568_clk;
wire [15:0] _U568_out;
wire [15:0] _U569_in;
wire _U569_clk;
wire [15:0] _U569_out;
wire [15:0] _U570_in;
wire _U570_clk;
wire [15:0] _U570_out;
wire [15:0] _U571_in;
wire _U571_clk;
wire [15:0] _U571_out;
wire [15:0] _U572_in;
wire [15:0] _U572_out;
wire [15:0] _U574_in;
wire _U574_clk;
wire [15:0] _U574_out;
wire [15:0] _U575_in;
wire _U575_clk;
wire [15:0] _U575_out;
wire [15:0] _U576_in;
wire _U576_clk;
wire [15:0] _U576_out;
wire [15:0] _U577_in;
wire _U577_clk;
wire [15:0] _U577_out;
wire [15:0] _U578_in;
wire _U578_clk;
wire [15:0] _U578_out;
wire [15:0] _U579_in;
wire [15:0] _U579_out;
wire [15:0] _U581_in;
wire _U581_clk;
wire [15:0] _U581_out;
wire [15:0] _U582_in;
wire _U582_clk;
wire [15:0] _U582_out;
wire [15:0] _U583_in;
wire _U583_clk;
wire [15:0] _U583_out;
wire [15:0] _U584_in;
wire _U584_clk;
wire [15:0] _U584_out;
wire [15:0] _U585_in;
wire _U585_clk;
wire [15:0] _U585_out;
wire [15:0] _U586_in;
wire _U586_clk;
wire [15:0] _U586_out;
wire [15:0] _U587_in;
wire [15:0] _U587_out;
wire [15:0] _U589_in;
wire _U589_clk;
wire [15:0] _U589_out;
wire [15:0] _U590_in;
wire _U590_clk;
wire [15:0] _U590_out;
wire [15:0] _U591_in;
wire _U591_clk;
wire [15:0] _U591_out;
wire [15:0] _U592_in;
wire _U592_clk;
wire [15:0] _U592_out;
wire [15:0] _U593_in;
wire _U593_clk;
wire [15:0] _U593_out;
wire [15:0] _U594_in;
wire _U594_clk;
wire [15:0] _U594_out;
wire [15:0] _U595_in;
wire [15:0] _U595_out;
wire [15:0] _U597_in;
wire _U597_clk;
wire [15:0] _U597_out;
wire [15:0] _U598_in;
wire _U598_clk;
wire [15:0] _U598_out;
wire [15:0] _U599_in;
wire _U599_clk;
wire [15:0] _U599_out;
wire [15:0] _U600_in;
wire _U600_clk;
wire [15:0] _U600_out;
wire [15:0] _U601_in;
wire _U601_clk;
wire [15:0] _U601_out;
wire [15:0] _U602_in;
wire _U602_clk;
wire [15:0] _U602_out;
wire [15:0] _U603_in;
wire _U603_clk;
wire [15:0] _U603_out;
wire [15:0] _U604_in;
wire [15:0] _U604_out;
wire [15:0] _U606_in;
wire _U606_clk;
wire [15:0] _U606_out;
wire [15:0] _U607_in;
wire _U607_clk;
wire [15:0] _U607_out;
wire [15:0] _U608_in;
wire _U608_clk;
wire [15:0] _U608_out;
wire [15:0] _U609_in;
wire _U609_clk;
wire [15:0] _U609_out;
wire [15:0] _U610_in;
wire _U610_clk;
wire [15:0] _U610_out;
wire [15:0] _U611_in;
wire _U611_clk;
wire [15:0] _U611_out;
wire [15:0] _U612_in;
wire _U612_clk;
wire [15:0] _U612_out;
assign _U412_in = _U428_out;
_U412_pt__U413 _U412 (
    .in(_U412_in),
    .out(_U412_out)
);
assign _U414_in = 16'(_U525_out * _U527_out);
assign _U414_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U414 (
    .in(_U414_in),
    .clk(_U414_clk),
    .out(_U414_out)
);
assign _U415_in = _U414_out;
assign _U415_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U415 (
    .in(_U415_in),
    .clk(_U415_clk),
    .out(_U415_out)
);
assign _U416_in = _U415_out;
assign _U416_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U416 (
    .in(_U416_in),
    .clk(_U416_clk),
    .out(_U416_out)
);
assign _U417_in = _U416_out;
assign _U417_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U417 (
    .in(_U417_in),
    .clk(_U417_clk),
    .out(_U417_out)
);
assign _U418_in = _U417_out;
assign _U418_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U418 (
    .in(_U418_in),
    .clk(_U418_clk),
    .out(_U418_out)
);
assign _U419_in = _U418_out;
assign _U419_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U419 (
    .in(_U419_in),
    .clk(_U419_clk),
    .out(_U419_out)
);
assign _U420_in = _U419_out;
assign _U420_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U420 (
    .in(_U420_in),
    .clk(_U420_clk),
    .out(_U420_out)
);
assign _U421_in = _U420_out;
assign _U421_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U421 (
    .in(_U421_in),
    .clk(_U421_clk),
    .out(_U421_out)
);
assign _U422_in = _U421_out;
assign _U422_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U422 (
    .in(_U422_in),
    .clk(_U422_clk),
    .out(_U422_out)
);
assign _U423_in = _U422_out;
assign _U423_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U423 (
    .in(_U423_in),
    .clk(_U423_clk),
    .out(_U423_out)
);
assign _U424_in = _U423_out;
assign _U424_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U424 (
    .in(_U424_in),
    .clk(_U424_clk),
    .out(_U424_out)
);
assign _U425_in = _U424_out;
assign _U425_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U425 (
    .in(_U425_in),
    .clk(_U425_clk),
    .out(_U425_out)
);
assign _U426_in = _U425_out;
assign _U426_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U426 (
    .in(_U426_in),
    .clk(_U426_clk),
    .out(_U426_out)
);
assign _U427_in = _U426_out;
assign _U427_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U427 (
    .in(_U427_in),
    .clk(_U427_clk),
    .out(_U427_out)
);
assign _U428_in = _U427_out;
assign _U428_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U428 (
    .in(_U428_in),
    .clk(_U428_clk),
    .out(_U428_out)
);
assign _U429_in = _U431_out;
_U429_pt__U430 _U429 (
    .in(_U429_in),
    .out(_U429_out)
);
assign _U431_in = 16'(_U509_out + _U451_out);
assign _U431_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U431 (
    .in(_U431_in),
    .clk(_U431_clk),
    .out(_U431_out)
);
assign _U432_in = 16'(_U412_out + _U429_out);
_U432_pt__U433 _U432 (
    .in(_U432_in),
    .out(out_conv_stencil)
);
assign _U434_in = _U447_out;
_U434_pt__U435 _U434 (
    .in(_U434_in),
    .out(_U434_out)
);
assign _U436_in = 16'(_U529_out * _U532_out);
assign _U436_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U436 (
    .in(_U436_in),
    .clk(_U436_clk),
    .out(_U436_out)
);
assign _U437_in = _U436_out;
assign _U437_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U437 (
    .in(_U437_in),
    .clk(_U437_clk),
    .out(_U437_out)
);
assign _U438_in = _U437_out;
assign _U438_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U438 (
    .in(_U438_in),
    .clk(_U438_clk),
    .out(_U438_out)
);
assign _U439_in = _U438_out;
assign _U439_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U439 (
    .in(_U439_in),
    .clk(_U439_clk),
    .out(_U439_out)
);
assign _U440_in = _U439_out;
assign _U440_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U440 (
    .in(_U440_in),
    .clk(_U440_clk),
    .out(_U440_out)
);
assign _U441_in = _U440_out;
assign _U441_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U441 (
    .in(_U441_in),
    .clk(_U441_clk),
    .out(_U441_out)
);
assign _U442_in = _U441_out;
assign _U442_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U442 (
    .in(_U442_in),
    .clk(_U442_clk),
    .out(_U442_out)
);
assign _U443_in = _U442_out;
assign _U443_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U443 (
    .in(_U443_in),
    .clk(_U443_clk),
    .out(_U443_out)
);
assign _U444_in = _U443_out;
assign _U444_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U444 (
    .in(_U444_in),
    .clk(_U444_clk),
    .out(_U444_out)
);
assign _U445_in = _U444_out;
assign _U445_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U445 (
    .in(_U445_in),
    .clk(_U445_clk),
    .out(_U445_out)
);
assign _U446_in = _U445_out;
assign _U446_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U446 (
    .in(_U446_in),
    .clk(_U446_clk),
    .out(_U446_out)
);
assign _U447_in = _U446_out;
assign _U447_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U447 (
    .in(_U447_in),
    .clk(_U447_clk),
    .out(_U447_out)
);
assign _U448_in = _U450_out;
_U448_pt__U449 _U448 (
    .in(_U448_in),
    .out(_U448_out)
);
assign _U450_in = 16'(_U454_out + _U466_out);
assign _U450_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U450 (
    .in(_U450_in),
    .clk(_U450_clk),
    .out(_U450_out)
);
assign _U451_in = _U453_out;
_U451_pt__U452 _U451 (
    .in(_U451_in),
    .out(_U451_out)
);
assign _U453_in = 16'(_U434_out + _U448_out);
assign _U453_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U453 (
    .in(_U453_in),
    .clk(_U453_clk),
    .out(_U453_out)
);
assign _U454_in = _U465_out;
_U454_pt__U455 _U454 (
    .in(_U454_in),
    .out(_U454_out)
);
assign _U456_in = 16'(_U535_out * _U539_out);
assign _U456_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U456 (
    .in(_U456_in),
    .clk(_U456_clk),
    .out(_U456_out)
);
assign _U457_in = _U456_out;
assign _U457_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U457 (
    .in(_U457_in),
    .clk(_U457_clk),
    .out(_U457_out)
);
assign _U458_in = _U457_out;
assign _U458_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U458 (
    .in(_U458_in),
    .clk(_U458_clk),
    .out(_U458_out)
);
assign _U459_in = _U458_out;
assign _U459_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U459 (
    .in(_U459_in),
    .clk(_U459_clk),
    .out(_U459_out)
);
assign _U460_in = _U459_out;
assign _U460_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U460 (
    .in(_U460_in),
    .clk(_U460_clk),
    .out(_U460_out)
);
assign _U461_in = _U460_out;
assign _U461_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U461 (
    .in(_U461_in),
    .clk(_U461_clk),
    .out(_U461_out)
);
assign _U462_in = _U461_out;
assign _U462_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U462 (
    .in(_U462_in),
    .clk(_U462_clk),
    .out(_U462_out)
);
assign _U463_in = _U462_out;
assign _U463_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U463 (
    .in(_U463_in),
    .clk(_U463_clk),
    .out(_U463_out)
);
assign _U464_in = _U463_out;
assign _U464_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U464 (
    .in(_U464_in),
    .clk(_U464_clk),
    .out(_U464_out)
);
assign _U465_in = _U464_out;
assign _U465_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U465 (
    .in(_U465_in),
    .clk(_U465_clk),
    .out(_U465_out)
);
assign _U466_in = _U468_out;
_U466_pt__U467 _U466 (
    .in(_U466_in),
    .out(_U466_out)
);
assign _U468_in = 16'(_U469_out + _U479_out);
assign _U468_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U468 (
    .in(_U468_in),
    .clk(_U468_clk),
    .out(_U468_out)
);
assign _U469_in = _U478_out;
_U469_pt__U470 _U469 (
    .in(_U469_in),
    .out(_U469_out)
);
assign _U471_in = 16'(_U543_out * _U548_out);
assign _U471_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U471 (
    .in(_U471_in),
    .clk(_U471_clk),
    .out(_U471_out)
);
assign _U472_in = _U471_out;
assign _U472_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U472 (
    .in(_U472_in),
    .clk(_U472_clk),
    .out(_U472_out)
);
assign _U473_in = _U472_out;
assign _U473_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U473 (
    .in(_U473_in),
    .clk(_U473_clk),
    .out(_U473_out)
);
assign _U474_in = _U473_out;
assign _U474_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U474 (
    .in(_U474_in),
    .clk(_U474_clk),
    .out(_U474_out)
);
assign _U475_in = _U474_out;
assign _U475_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U475 (
    .in(_U475_in),
    .clk(_U475_clk),
    .out(_U475_out)
);
assign _U476_in = _U475_out;
assign _U476_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U476 (
    .in(_U476_in),
    .clk(_U476_clk),
    .out(_U476_out)
);
assign _U477_in = _U476_out;
assign _U477_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U477 (
    .in(_U477_in),
    .clk(_U477_clk),
    .out(_U477_out)
);
assign _U478_in = _U477_out;
assign _U478_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U478 (
    .in(_U478_in),
    .clk(_U478_clk),
    .out(_U478_out)
);
assign _U479_in = _U481_out;
_U479_pt__U480 _U479 (
    .in(_U479_in),
    .out(_U479_out)
);
assign _U481_in = 16'(_U482_out + _U490_out);
assign _U481_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U481 (
    .in(_U481_in),
    .clk(_U481_clk),
    .out(_U481_out)
);
assign _U482_in = _U489_out;
_U482_pt__U483 _U482 (
    .in(_U482_in),
    .out(_U482_out)
);
assign _U484_in = 16'(_U553_out * _U559_out);
assign _U484_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U484 (
    .in(_U484_in),
    .clk(_U484_clk),
    .out(_U484_out)
);
assign _U485_in = _U484_out;
assign _U485_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U485 (
    .in(_U485_in),
    .clk(_U485_clk),
    .out(_U485_out)
);
assign _U486_in = _U485_out;
assign _U486_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U486 (
    .in(_U486_in),
    .clk(_U486_clk),
    .out(_U486_out)
);
assign _U487_in = _U486_out;
assign _U487_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U487 (
    .in(_U487_in),
    .clk(_U487_clk),
    .out(_U487_out)
);
assign _U488_in = _U487_out;
assign _U488_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U488 (
    .in(_U488_in),
    .clk(_U488_clk),
    .out(_U488_out)
);
assign _U489_in = _U488_out;
assign _U489_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U489 (
    .in(_U489_in),
    .clk(_U489_clk),
    .out(_U489_out)
);
assign _U490_in = _U492_out;
_U490_pt__U491 _U490 (
    .in(_U490_in),
    .out(_U490_out)
);
assign _U492_in = 16'(_U493_out + _U499_out);
assign _U492_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U492 (
    .in(_U492_in),
    .clk(_U492_clk),
    .out(_U492_out)
);
assign _U493_in = _U498_out;
_U493_pt__U494 _U493 (
    .in(_U493_in),
    .out(_U493_out)
);
assign _U495_in = 16'(_U565_out * _U572_out);
assign _U495_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U495 (
    .in(_U495_in),
    .clk(_U495_clk),
    .out(_U495_out)
);
assign _U496_in = _U495_out;
assign _U496_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U496 (
    .in(_U496_in),
    .clk(_U496_clk),
    .out(_U496_out)
);
assign _U497_in = _U496_out;
assign _U497_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U497 (
    .in(_U497_in),
    .clk(_U497_clk),
    .out(_U497_out)
);
assign _U498_in = _U497_out;
assign _U498_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U498 (
    .in(_U498_in),
    .clk(_U498_clk),
    .out(_U498_out)
);
assign _U499_in = _U501_out;
_U499_pt__U500 _U499 (
    .in(_U499_in),
    .out(_U499_out)
);
assign _U501_in = 16'(_U502_out + _U506_out);
assign _U501_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U501 (
    .in(_U501_in),
    .clk(_U501_clk),
    .out(_U501_out)
);
assign _U502_in = _U505_out;
_U502_pt__U503 _U502 (
    .in(_U502_in),
    .out(_U502_out)
);
assign _U504_in = 16'(_U579_out * _U587_out);
assign _U504_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U504 (
    .in(_U504_in),
    .clk(_U504_clk),
    .out(_U504_out)
);
assign _U505_in = _U504_out;
assign _U505_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U505 (
    .in(_U505_in),
    .clk(_U505_clk),
    .out(_U505_out)
);
assign _U506_in = _U508_out;
_U506_pt__U507 _U506 (
    .in(_U506_in),
    .out(_U506_out)
);
assign _U508_in = 16'(_U595_out * _U604_out);
assign _U508_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U508 (
    .in(_U508_in),
    .clk(_U508_clk),
    .out(_U508_out)
);
assign _U509_in = _U524_out;
_U509_pt__U510 _U509 (
    .in(_U509_in),
    .out(_U509_out)
);
assign _U511_in = in0_conv_stencil[0];
assign _U511_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U511 (
    .in(_U511_in),
    .clk(_U511_clk),
    .out(_U511_out)
);
assign _U512_in = _U511_out;
assign _U512_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U512 (
    .in(_U512_in),
    .clk(_U512_clk),
    .out(_U512_out)
);
assign _U513_in = _U512_out;
assign _U513_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U513 (
    .in(_U513_in),
    .clk(_U513_clk),
    .out(_U513_out)
);
assign _U514_in = _U513_out;
assign _U514_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U514 (
    .in(_U514_in),
    .clk(_U514_clk),
    .out(_U514_out)
);
assign _U515_in = _U514_out;
assign _U515_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U515 (
    .in(_U515_in),
    .clk(_U515_clk),
    .out(_U515_out)
);
assign _U516_in = _U515_out;
assign _U516_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U516 (
    .in(_U516_in),
    .clk(_U516_clk),
    .out(_U516_out)
);
assign _U517_in = _U516_out;
assign _U517_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U517 (
    .in(_U517_in),
    .clk(_U517_clk),
    .out(_U517_out)
);
assign _U518_in = _U517_out;
assign _U518_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U518 (
    .in(_U518_in),
    .clk(_U518_clk),
    .out(_U518_out)
);
assign _U519_in = _U518_out;
assign _U519_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U519 (
    .in(_U519_in),
    .clk(_U519_clk),
    .out(_U519_out)
);
assign _U520_in = _U519_out;
assign _U520_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U520 (
    .in(_U520_in),
    .clk(_U520_clk),
    .out(_U520_out)
);
assign _U521_in = _U520_out;
assign _U521_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U521 (
    .in(_U521_in),
    .clk(_U521_clk),
    .out(_U521_out)
);
assign _U522_in = _U521_out;
assign _U522_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U522 (
    .in(_U522_in),
    .clk(_U522_clk),
    .out(_U522_out)
);
assign _U523_in = _U522_out;
assign _U523_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U523 (
    .in(_U523_in),
    .clk(_U523_clk),
    .out(_U523_out)
);
assign _U524_in = _U523_out;
assign _U524_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U524 (
    .in(_U524_in),
    .clk(_U524_clk),
    .out(_U524_out)
);
assign _U525_in = in2_hw_kernel_global_wrapper_stencil[0];
_U525_pt__U526 _U525 (
    .in(_U525_in),
    .out(_U525_out)
);
assign _U527_in = in1_hw_input_global_wrapper_stencil[0];
_U527_pt__U528 _U527 (
    .in(_U527_in),
    .out(_U527_out)
);
assign _U529_in = _U531_out;
_U529_pt__U530 _U529 (
    .in(_U529_in),
    .out(_U529_out)
);
assign _U531_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U531_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U531 (
    .in(_U531_in),
    .clk(_U531_clk),
    .out(_U531_out)
);
assign _U532_in = _U534_out;
_U532_pt__U533 _U532 (
    .in(_U532_in),
    .out(_U532_out)
);
assign _U534_in = in1_hw_input_global_wrapper_stencil[1];
assign _U534_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U534 (
    .in(_U534_in),
    .clk(_U534_clk),
    .out(_U534_out)
);
assign _U535_in = _U538_out;
_U535_pt__U536 _U535 (
    .in(_U535_in),
    .out(_U535_out)
);
assign _U537_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U537_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U537 (
    .in(_U537_in),
    .clk(_U537_clk),
    .out(_U537_out)
);
assign _U538_in = _U537_out;
assign _U538_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U538 (
    .in(_U538_in),
    .clk(_U538_clk),
    .out(_U538_out)
);
assign _U539_in = _U542_out;
_U539_pt__U540 _U539 (
    .in(_U539_in),
    .out(_U539_out)
);
assign _U541_in = in1_hw_input_global_wrapper_stencil[2];
assign _U541_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U541 (
    .in(_U541_in),
    .clk(_U541_clk),
    .out(_U541_out)
);
assign _U542_in = _U541_out;
assign _U542_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U542 (
    .in(_U542_in),
    .clk(_U542_clk),
    .out(_U542_out)
);
assign _U543_in = _U547_out;
_U543_pt__U544 _U543 (
    .in(_U543_in),
    .out(_U543_out)
);
assign _U545_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U545_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U545 (
    .in(_U545_in),
    .clk(_U545_clk),
    .out(_U545_out)
);
assign _U546_in = _U545_out;
assign _U546_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U546 (
    .in(_U546_in),
    .clk(_U546_clk),
    .out(_U546_out)
);
assign _U547_in = _U546_out;
assign _U547_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U547 (
    .in(_U547_in),
    .clk(_U547_clk),
    .out(_U547_out)
);
assign _U548_in = _U552_out;
_U548_pt__U549 _U548 (
    .in(_U548_in),
    .out(_U548_out)
);
assign _U550_in = in1_hw_input_global_wrapper_stencil[3];
assign _U550_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U550 (
    .in(_U550_in),
    .clk(_U550_clk),
    .out(_U550_out)
);
assign _U551_in = _U550_out;
assign _U551_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U551 (
    .in(_U551_in),
    .clk(_U551_clk),
    .out(_U551_out)
);
assign _U552_in = _U551_out;
assign _U552_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U552 (
    .in(_U552_in),
    .clk(_U552_clk),
    .out(_U552_out)
);
assign _U553_in = _U558_out;
_U553_pt__U554 _U553 (
    .in(_U553_in),
    .out(_U553_out)
);
assign _U555_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U555_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U555 (
    .in(_U555_in),
    .clk(_U555_clk),
    .out(_U555_out)
);
assign _U556_in = _U555_out;
assign _U556_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U556 (
    .in(_U556_in),
    .clk(_U556_clk),
    .out(_U556_out)
);
assign _U557_in = _U556_out;
assign _U557_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U557 (
    .in(_U557_in),
    .clk(_U557_clk),
    .out(_U557_out)
);
assign _U558_in = _U557_out;
assign _U558_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U558 (
    .in(_U558_in),
    .clk(_U558_clk),
    .out(_U558_out)
);
assign _U559_in = _U564_out;
_U559_pt__U560 _U559 (
    .in(_U559_in),
    .out(_U559_out)
);
assign _U561_in = in1_hw_input_global_wrapper_stencil[4];
assign _U561_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U561 (
    .in(_U561_in),
    .clk(_U561_clk),
    .out(_U561_out)
);
assign _U562_in = _U561_out;
assign _U562_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U562 (
    .in(_U562_in),
    .clk(_U562_clk),
    .out(_U562_out)
);
assign _U563_in = _U562_out;
assign _U563_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U563 (
    .in(_U563_in),
    .clk(_U563_clk),
    .out(_U563_out)
);
assign _U564_in = _U563_out;
assign _U564_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U564 (
    .in(_U564_in),
    .clk(_U564_clk),
    .out(_U564_out)
);
assign _U565_in = _U571_out;
_U565_pt__U566 _U565 (
    .in(_U565_in),
    .out(_U565_out)
);
assign _U567_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U567_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U567 (
    .in(_U567_in),
    .clk(_U567_clk),
    .out(_U567_out)
);
assign _U568_in = _U567_out;
assign _U568_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U568 (
    .in(_U568_in),
    .clk(_U568_clk),
    .out(_U568_out)
);
assign _U569_in = _U568_out;
assign _U569_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U569 (
    .in(_U569_in),
    .clk(_U569_clk),
    .out(_U569_out)
);
assign _U570_in = _U569_out;
assign _U570_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U570 (
    .in(_U570_in),
    .clk(_U570_clk),
    .out(_U570_out)
);
assign _U571_in = _U570_out;
assign _U571_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U571 (
    .in(_U571_in),
    .clk(_U571_clk),
    .out(_U571_out)
);
assign _U572_in = _U578_out;
_U572_pt__U573 _U572 (
    .in(_U572_in),
    .out(_U572_out)
);
assign _U574_in = in1_hw_input_global_wrapper_stencil[5];
assign _U574_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U574 (
    .in(_U574_in),
    .clk(_U574_clk),
    .out(_U574_out)
);
assign _U575_in = _U574_out;
assign _U575_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U575 (
    .in(_U575_in),
    .clk(_U575_clk),
    .out(_U575_out)
);
assign _U576_in = _U575_out;
assign _U576_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U576 (
    .in(_U576_in),
    .clk(_U576_clk),
    .out(_U576_out)
);
assign _U577_in = _U576_out;
assign _U577_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U577 (
    .in(_U577_in),
    .clk(_U577_clk),
    .out(_U577_out)
);
assign _U578_in = _U577_out;
assign _U578_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U578 (
    .in(_U578_in),
    .clk(_U578_clk),
    .out(_U578_out)
);
assign _U579_in = _U586_out;
_U579_pt__U580 _U579 (
    .in(_U579_in),
    .out(_U579_out)
);
assign _U581_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U581_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U581 (
    .in(_U581_in),
    .clk(_U581_clk),
    .out(_U581_out)
);
assign _U582_in = _U581_out;
assign _U582_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U582 (
    .in(_U582_in),
    .clk(_U582_clk),
    .out(_U582_out)
);
assign _U583_in = _U582_out;
assign _U583_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U583 (
    .in(_U583_in),
    .clk(_U583_clk),
    .out(_U583_out)
);
assign _U584_in = _U583_out;
assign _U584_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U584 (
    .in(_U584_in),
    .clk(_U584_clk),
    .out(_U584_out)
);
assign _U585_in = _U584_out;
assign _U585_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U585 (
    .in(_U585_in),
    .clk(_U585_clk),
    .out(_U585_out)
);
assign _U586_in = _U585_out;
assign _U586_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U586 (
    .in(_U586_in),
    .clk(_U586_clk),
    .out(_U586_out)
);
assign _U587_in = _U594_out;
_U587_pt__U588 _U587 (
    .in(_U587_in),
    .out(_U587_out)
);
assign _U589_in = in1_hw_input_global_wrapper_stencil[6];
assign _U589_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U589 (
    .in(_U589_in),
    .clk(_U589_clk),
    .out(_U589_out)
);
assign _U590_in = _U589_out;
assign _U590_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U590 (
    .in(_U590_in),
    .clk(_U590_clk),
    .out(_U590_out)
);
assign _U591_in = _U590_out;
assign _U591_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U591 (
    .in(_U591_in),
    .clk(_U591_clk),
    .out(_U591_out)
);
assign _U592_in = _U591_out;
assign _U592_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U592 (
    .in(_U592_in),
    .clk(_U592_clk),
    .out(_U592_out)
);
assign _U593_in = _U592_out;
assign _U593_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U593 (
    .in(_U593_in),
    .clk(_U593_clk),
    .out(_U593_out)
);
assign _U594_in = _U593_out;
assign _U594_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U594 (
    .in(_U594_in),
    .clk(_U594_clk),
    .out(_U594_out)
);
assign _U595_in = _U603_out;
_U595_pt__U596 _U595 (
    .in(_U595_in),
    .out(_U595_out)
);
assign _U597_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U597_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U597 (
    .in(_U597_in),
    .clk(_U597_clk),
    .out(_U597_out)
);
assign _U598_in = _U597_out;
assign _U598_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U598 (
    .in(_U598_in),
    .clk(_U598_clk),
    .out(_U598_out)
);
assign _U599_in = _U598_out;
assign _U599_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U599 (
    .in(_U599_in),
    .clk(_U599_clk),
    .out(_U599_out)
);
assign _U600_in = _U599_out;
assign _U600_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U600 (
    .in(_U600_in),
    .clk(_U600_clk),
    .out(_U600_out)
);
assign _U601_in = _U600_out;
assign _U601_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U601 (
    .in(_U601_in),
    .clk(_U601_clk),
    .out(_U601_out)
);
assign _U602_in = _U601_out;
assign _U602_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U602 (
    .in(_U602_in),
    .clk(_U602_clk),
    .out(_U602_out)
);
assign _U603_in = _U602_out;
assign _U603_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U603 (
    .in(_U603_in),
    .clk(_U603_clk),
    .out(_U603_out)
);
assign _U604_in = _U612_out;
_U604_pt__U605 _U604 (
    .in(_U604_in),
    .out(_U604_out)
);
assign _U606_in = in1_hw_input_global_wrapper_stencil[7];
assign _U606_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U606 (
    .in(_U606_in),
    .clk(_U606_clk),
    .out(_U606_out)
);
assign _U607_in = _U606_out;
assign _U607_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U607 (
    .in(_U607_in),
    .clk(_U607_clk),
    .out(_U607_out)
);
assign _U608_in = _U607_out;
assign _U608_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U608 (
    .in(_U608_in),
    .clk(_U608_clk),
    .out(_U608_out)
);
assign _U609_in = _U608_out;
assign _U609_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U609 (
    .in(_U609_in),
    .clk(_U609_clk),
    .out(_U609_out)
);
assign _U610_in = _U609_out;
assign _U610_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U610 (
    .in(_U610_in),
    .clk(_U610_clk),
    .out(_U610_out)
);
assign _U611_in = _U610_out;
assign _U611_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U611 (
    .in(_U611_in),
    .clk(_U611_clk),
    .out(_U611_out)
);
assign _U612_in = _U611_out;
assign _U612_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U612 (
    .in(_U612_in),
    .clk(_U612_clk),
    .out(_U612_out)
);
endmodule

module cu_op_hcompute_conv_stencil_3 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
hcompute_conv_stencil_3_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U396_pt__U397 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U393_pt__U394 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U388_pt__U389 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U381_pt__U382 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U378_pt__U379 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U364_pt__U365 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U362_pt__U363 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U359_pt__U360 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U357_pt__U358 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U353_pt__U354 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U348_pt__U349 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U337_pt__U338 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U334_pt__U335 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U331_pt__U332 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U328_pt__U329 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U323_pt__U324 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U317_pt__U318 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U313_pt__U314 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U303_pt__U304 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U2_pt__U3 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_1_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U2_in;
assign _U2_in = 16'h0000;
_U2_pt__U3 _U2 (
    .in(_U2_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil_1 (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_1_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U292_pt__U293 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U282_pt__U283 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U280_pt__U281 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U27_pt__U28 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U274_pt__U275 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U268_pt__U269 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U256_pt__U257 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U252_pt__U253 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U244_pt__U245 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U241_pt__U242 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U238_pt__U239 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U235_pt__U236 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U228_pt__U229 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U223_pt__U224 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U211_pt__U212 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_4_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U211_in;
wire [15:0] _U211_out;
wire [15:0] _U213_in;
wire _U213_clk;
wire [15:0] _U213_out;
wire [15:0] _U214_in;
wire _U214_clk;
wire [15:0] _U214_out;
wire [15:0] _U215_in;
wire _U215_clk;
wire [15:0] _U215_out;
wire [15:0] _U216_in;
wire _U216_clk;
wire [15:0] _U216_out;
wire [15:0] _U217_in;
wire _U217_clk;
wire [15:0] _U217_out;
wire [15:0] _U218_in;
wire _U218_clk;
wire [15:0] _U218_out;
wire [15:0] _U219_in;
wire _U219_clk;
wire [15:0] _U219_out;
wire [15:0] _U220_in;
wire _U220_clk;
wire [15:0] _U220_out;
wire [15:0] _U221_in;
wire _U221_clk;
wire [15:0] _U221_out;
wire [15:0] _U222_in;
wire _U222_clk;
wire [15:0] _U222_out;
wire [15:0] _U223_in;
wire [15:0] _U223_out;
wire [15:0] _U225_in;
wire _U225_clk;
wire [15:0] _U225_out;
wire [15:0] _U226_in;
wire _U226_clk;
wire [15:0] _U226_out;
wire [15:0] _U227_in;
wire _U227_clk;
wire [15:0] _U227_out;
wire [15:0] _U228_in;
wire [15:0] _U228_out;
wire [15:0] _U230_in;
wire _U230_clk;
wire [15:0] _U230_out;
wire [15:0] _U231_in;
wire _U231_clk;
wire [15:0] _U231_out;
wire [15:0] _U232_in;
wire _U232_clk;
wire [15:0] _U232_out;
wire [15:0] _U233_in;
wire _U233_clk;
wire [15:0] _U233_out;
wire [15:0] _U234_in;
wire _U234_clk;
wire [15:0] _U234_out;
wire [15:0] _U235_in;
wire [15:0] _U235_out;
wire [15:0] _U237_in;
wire _U237_clk;
wire [15:0] _U237_out;
wire [15:0] _U238_in;
wire [15:0] _U238_out;
wire [15:0] _U240_in;
wire _U240_clk;
wire [15:0] _U240_out;
wire [15:0] _U241_in;
wire [15:0] _U241_out;
wire [15:0] _U243_in;
wire _U243_clk;
wire [15:0] _U243_out;
wire [15:0] _U244_in;
wire [15:0] _U244_out;
wire [15:0] _U246_in;
wire _U246_clk;
wire [15:0] _U246_out;
wire [15:0] _U247_in;
wire _U247_clk;
wire [15:0] _U247_out;
wire [15:0] _U248_in;
wire _U248_clk;
wire [15:0] _U248_out;
wire [15:0] _U249_in;
wire _U249_clk;
wire [15:0] _U249_out;
wire [15:0] _U250_in;
wire _U250_clk;
wire [15:0] _U250_out;
wire [15:0] _U251_in;
wire _U251_clk;
wire [15:0] _U251_out;
wire [15:0] _U252_in;
wire [15:0] _U252_out;
wire [15:0] _U254_in;
wire _U254_clk;
wire [15:0] _U254_out;
wire [15:0] _U255_in;
wire _U255_clk;
wire [15:0] _U255_out;
wire [15:0] _U256_in;
wire [15:0] _U256_out;
wire [15:0] _U258_in;
wire _U258_clk;
wire [15:0] _U258_out;
wire [15:0] _U259_in;
wire _U259_clk;
wire [15:0] _U259_out;
wire [15:0] _U260_in;
wire _U260_clk;
wire [15:0] _U260_out;
wire [15:0] _U261_in;
wire _U261_clk;
wire [15:0] _U261_out;
wire [15:0] _U262_in;
wire _U262_clk;
wire [15:0] _U262_out;
wire [15:0] _U263_in;
wire _U263_clk;
wire [15:0] _U263_out;
wire [15:0] _U264_in;
wire _U264_clk;
wire [15:0] _U264_out;
wire [15:0] _U265_in;
wire _U265_clk;
wire [15:0] _U265_out;
wire [15:0] _U266_in;
wire _U266_clk;
wire [15:0] _U266_out;
wire [15:0] _U267_in;
wire _U267_clk;
wire [15:0] _U267_out;
wire [15:0] _U268_in;
wire [15:0] _U268_out;
wire [15:0] _U270_in;
wire _U270_clk;
wire [15:0] _U270_out;
wire [15:0] _U271_in;
wire _U271_clk;
wire [15:0] _U271_out;
wire [15:0] _U272_in;
wire _U272_clk;
wire [15:0] _U272_out;
wire [15:0] _U273_in;
wire _U273_clk;
wire [15:0] _U273_out;
wire [15:0] _U274_in;
wire [15:0] _U274_out;
wire [15:0] _U276_in;
wire _U276_clk;
wire [15:0] _U276_out;
wire [15:0] _U277_in;
wire _U277_clk;
wire [15:0] _U277_out;
wire [15:0] _U278_in;
wire _U278_clk;
wire [15:0] _U278_out;
wire [15:0] _U279_in;
wire _U279_clk;
wire [15:0] _U279_out;
wire [15:0] _U280_in;
wire [15:0] _U282_in;
wire [15:0] _U282_out;
wire [15:0] _U284_in;
wire _U284_clk;
wire [15:0] _U284_out;
wire [15:0] _U285_in;
wire _U285_clk;
wire [15:0] _U285_out;
wire [15:0] _U286_in;
wire _U286_clk;
wire [15:0] _U286_out;
wire [15:0] _U287_in;
wire _U287_clk;
wire [15:0] _U287_out;
wire [15:0] _U288_in;
wire _U288_clk;
wire [15:0] _U288_out;
wire [15:0] _U289_in;
wire _U289_clk;
wire [15:0] _U289_out;
wire [15:0] _U290_in;
wire _U290_clk;
wire [15:0] _U290_out;
wire [15:0] _U291_in;
wire _U291_clk;
wire [15:0] _U291_out;
wire [15:0] _U292_in;
wire [15:0] _U292_out;
wire [15:0] _U294_in;
wire _U294_clk;
wire [15:0] _U294_out;
wire [15:0] _U295_in;
wire _U295_clk;
wire [15:0] _U295_out;
wire [15:0] _U296_in;
wire _U296_clk;
wire [15:0] _U296_out;
wire [15:0] _U297_in;
wire _U297_clk;
wire [15:0] _U297_out;
wire [15:0] _U298_in;
wire _U298_clk;
wire [15:0] _U298_out;
wire [15:0] _U299_in;
wire _U299_clk;
wire [15:0] _U299_out;
wire [15:0] _U300_in;
wire _U300_clk;
wire [15:0] _U300_out;
wire [15:0] _U301_in;
wire _U301_clk;
wire [15:0] _U301_out;
wire [15:0] _U302_in;
wire _U302_clk;
wire [15:0] _U302_out;
wire [15:0] _U303_in;
wire [15:0] _U303_out;
wire [15:0] _U305_in;
wire _U305_clk;
wire [15:0] _U305_out;
wire [15:0] _U306_in;
wire _U306_clk;
wire [15:0] _U306_out;
wire [15:0] _U307_in;
wire _U307_clk;
wire [15:0] _U307_out;
wire [15:0] _U308_in;
wire _U308_clk;
wire [15:0] _U308_out;
wire [15:0] _U309_in;
wire _U309_clk;
wire [15:0] _U309_out;
wire [15:0] _U310_in;
wire _U310_clk;
wire [15:0] _U310_out;
wire [15:0] _U311_in;
wire _U311_clk;
wire [15:0] _U311_out;
wire [15:0] _U312_in;
wire _U312_clk;
wire [15:0] _U312_out;
wire [15:0] _U313_in;
wire [15:0] _U313_out;
wire [15:0] _U315_in;
wire _U315_clk;
wire [15:0] _U315_out;
wire [15:0] _U316_in;
wire _U316_clk;
wire [15:0] _U316_out;
wire [15:0] _U317_in;
wire [15:0] _U317_out;
wire [15:0] _U319_in;
wire _U319_clk;
wire [15:0] _U319_out;
wire [15:0] _U320_in;
wire _U320_clk;
wire [15:0] _U320_out;
wire [15:0] _U321_in;
wire _U321_clk;
wire [15:0] _U321_out;
wire [15:0] _U322_in;
wire _U322_clk;
wire [15:0] _U322_out;
wire [15:0] _U323_in;
wire [15:0] _U323_out;
wire [15:0] _U325_in;
wire _U325_clk;
wire [15:0] _U325_out;
wire [15:0] _U326_in;
wire _U326_clk;
wire [15:0] _U326_out;
wire [15:0] _U327_in;
wire _U327_clk;
wire [15:0] _U327_out;
wire [15:0] _U328_in;
wire [15:0] _U328_out;
wire [15:0] _U330_in;
wire _U330_clk;
wire [15:0] _U330_out;
wire [15:0] _U331_in;
wire [15:0] _U331_out;
wire [15:0] _U333_in;
wire _U333_clk;
wire [15:0] _U333_out;
wire [15:0] _U334_in;
wire [15:0] _U334_out;
wire [15:0] _U336_in;
wire _U336_clk;
wire [15:0] _U336_out;
wire [15:0] _U337_in;
wire [15:0] _U337_out;
wire [15:0] _U339_in;
wire _U339_clk;
wire [15:0] _U339_out;
wire [15:0] _U340_in;
wire _U340_clk;
wire [15:0] _U340_out;
wire [15:0] _U341_in;
wire _U341_clk;
wire [15:0] _U341_out;
wire [15:0] _U342_in;
wire _U342_clk;
wire [15:0] _U342_out;
wire [15:0] _U343_in;
wire _U343_clk;
wire [15:0] _U343_out;
wire [15:0] _U344_in;
wire _U344_clk;
wire [15:0] _U344_out;
wire [15:0] _U345_in;
wire _U345_clk;
wire [15:0] _U345_out;
wire [15:0] _U346_in;
wire _U346_clk;
wire [15:0] _U346_out;
wire [15:0] _U347_in;
wire _U347_clk;
wire [15:0] _U347_out;
wire [15:0] _U348_in;
wire [15:0] _U348_out;
wire [15:0] _U350_in;
wire _U350_clk;
wire [15:0] _U350_out;
wire [15:0] _U351_in;
wire _U351_clk;
wire [15:0] _U351_out;
wire [15:0] _U352_in;
wire _U352_clk;
wire [15:0] _U352_out;
wire [15:0] _U353_in;
wire [15:0] _U353_out;
wire [15:0] _U355_in;
wire _U355_clk;
wire [15:0] _U355_out;
wire [15:0] _U356_in;
wire _U356_clk;
wire [15:0] _U356_out;
wire [15:0] _U357_in;
wire [15:0] _U357_out;
wire [15:0] _U359_in;
wire [15:0] _U359_out;
wire [15:0] _U361_in;
wire _U361_clk;
wire [15:0] _U361_out;
wire [15:0] _U362_in;
wire [15:0] _U362_out;
wire [15:0] _U364_in;
wire [15:0] _U364_out;
wire [15:0] _U366_in;
wire _U366_clk;
wire [15:0] _U366_out;
wire [15:0] _U367_in;
wire _U367_clk;
wire [15:0] _U367_out;
wire [15:0] _U368_in;
wire _U368_clk;
wire [15:0] _U368_out;
wire [15:0] _U369_in;
wire _U369_clk;
wire [15:0] _U369_out;
wire [15:0] _U370_in;
wire _U370_clk;
wire [15:0] _U370_out;
wire [15:0] _U371_in;
wire _U371_clk;
wire [15:0] _U371_out;
wire [15:0] _U372_in;
wire _U372_clk;
wire [15:0] _U372_out;
wire [15:0] _U373_in;
wire _U373_clk;
wire [15:0] _U373_out;
wire [15:0] _U374_in;
wire _U374_clk;
wire [15:0] _U374_out;
wire [15:0] _U375_in;
wire _U375_clk;
wire [15:0] _U375_out;
wire [15:0] _U376_in;
wire _U376_clk;
wire [15:0] _U376_out;
wire [15:0] _U377_in;
wire _U377_clk;
wire [15:0] _U377_out;
wire [15:0] _U378_in;
wire [15:0] _U378_out;
wire [15:0] _U380_in;
wire _U380_clk;
wire [15:0] _U380_out;
wire [15:0] _U381_in;
wire [15:0] _U381_out;
wire [15:0] _U383_in;
wire _U383_clk;
wire [15:0] _U383_out;
wire [15:0] _U384_in;
wire _U384_clk;
wire [15:0] _U384_out;
wire [15:0] _U385_in;
wire _U385_clk;
wire [15:0] _U385_out;
wire [15:0] _U386_in;
wire _U386_clk;
wire [15:0] _U386_out;
wire [15:0] _U387_in;
wire _U387_clk;
wire [15:0] _U387_out;
wire [15:0] _U388_in;
wire [15:0] _U388_out;
wire [15:0] _U390_in;
wire _U390_clk;
wire [15:0] _U390_out;
wire [15:0] _U391_in;
wire _U391_clk;
wire [15:0] _U391_out;
wire [15:0] _U392_in;
wire _U392_clk;
wire [15:0] _U392_out;
wire [15:0] _U393_in;
wire [15:0] _U393_out;
wire [15:0] _U395_in;
wire _U395_clk;
wire [15:0] _U395_out;
wire [15:0] _U396_in;
wire [15:0] _U396_out;
wire [15:0] _U398_in;
wire _U398_clk;
wire [15:0] _U398_out;
wire [15:0] _U399_in;
wire _U399_clk;
wire [15:0] _U399_out;
wire [15:0] _U400_in;
wire _U400_clk;
wire [15:0] _U400_out;
wire [15:0] _U401_in;
wire _U401_clk;
wire [15:0] _U401_out;
wire [15:0] _U402_in;
wire _U402_clk;
wire [15:0] _U402_out;
wire [15:0] _U403_in;
wire _U403_clk;
wire [15:0] _U403_out;
wire [15:0] _U404_in;
wire _U404_clk;
wire [15:0] _U404_out;
wire [15:0] _U405_in;
wire _U405_clk;
wire [15:0] _U405_out;
wire [15:0] _U406_in;
wire _U406_clk;
wire [15:0] _U406_out;
wire [15:0] _U407_in;
wire _U407_clk;
wire [15:0] _U407_out;
wire [15:0] _U408_in;
wire _U408_clk;
wire [15:0] _U408_out;
wire [15:0] _U409_in;
wire _U409_clk;
wire [15:0] _U409_out;
wire [15:0] _U410_in;
wire _U410_clk;
wire [15:0] _U410_out;
wire [15:0] _U411_in;
wire _U411_clk;
wire [15:0] _U411_out;
assign _U211_in = _U222_out;
_U211_pt__U212 _U211 (
    .in(_U211_in),
    .out(_U211_out)
);
assign _U213_in = in1_hw_input_global_wrapper_stencil[2];
assign _U213_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U213 (
    .in(_U213_in),
    .clk(_U213_clk),
    .out(_U213_out)
);
assign _U214_in = _U213_out;
assign _U214_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U214 (
    .in(_U214_in),
    .clk(_U214_clk),
    .out(_U214_out)
);
assign _U215_in = _U214_out;
assign _U215_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U215 (
    .in(_U215_in),
    .clk(_U215_clk),
    .out(_U215_out)
);
assign _U216_in = _U215_out;
assign _U216_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U216 (
    .in(_U216_in),
    .clk(_U216_clk),
    .out(_U216_out)
);
assign _U217_in = _U216_out;
assign _U217_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U217 (
    .in(_U217_in),
    .clk(_U217_clk),
    .out(_U217_out)
);
assign _U218_in = _U217_out;
assign _U218_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U218 (
    .in(_U218_in),
    .clk(_U218_clk),
    .out(_U218_out)
);
assign _U219_in = _U218_out;
assign _U219_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U219 (
    .in(_U219_in),
    .clk(_U219_clk),
    .out(_U219_out)
);
assign _U220_in = _U219_out;
assign _U220_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U220 (
    .in(_U220_in),
    .clk(_U220_clk),
    .out(_U220_out)
);
assign _U221_in = _U220_out;
assign _U221_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U221 (
    .in(_U221_in),
    .clk(_U221_clk),
    .out(_U221_out)
);
assign _U222_in = _U221_out;
assign _U222_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U222 (
    .in(_U222_in),
    .clk(_U222_clk),
    .out(_U222_out)
);
assign _U223_in = _U227_out;
_U223_pt__U224 _U223 (
    .in(_U223_in),
    .out(_U223_out)
);
assign _U225_in = in1_hw_input_global_wrapper_stencil[7];
assign _U225_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U225 (
    .in(_U225_in),
    .clk(_U225_clk),
    .out(_U225_out)
);
assign _U226_in = _U225_out;
assign _U226_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U226 (
    .in(_U226_in),
    .clk(_U226_clk),
    .out(_U226_out)
);
assign _U227_in = _U226_out;
assign _U227_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U227 (
    .in(_U227_in),
    .clk(_U227_clk),
    .out(_U227_out)
);
assign _U228_in = _U234_out;
_U228_pt__U229 _U228 (
    .in(_U228_in),
    .out(_U228_out)
);
assign _U230_in = 16'(_U282_out * _U303_out);
assign _U230_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U230 (
    .in(_U230_in),
    .clk(_U230_clk),
    .out(_U230_out)
);
assign _U231_in = _U230_out;
assign _U231_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U231 (
    .in(_U231_in),
    .clk(_U231_clk),
    .out(_U231_out)
);
assign _U232_in = _U231_out;
assign _U232_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U232 (
    .in(_U232_in),
    .clk(_U232_clk),
    .out(_U232_out)
);
assign _U233_in = _U232_out;
assign _U233_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U233 (
    .in(_U233_in),
    .clk(_U233_clk),
    .out(_U233_out)
);
assign _U234_in = _U233_out;
assign _U234_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U234 (
    .in(_U234_in),
    .clk(_U234_clk),
    .out(_U234_out)
);
assign _U235_in = _U237_out;
_U235_pt__U236 _U235 (
    .in(_U235_in),
    .out(_U235_out)
);
assign _U237_in = 16'(_U256_out * _U211_out);
assign _U237_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U237 (
    .in(_U237_in),
    .clk(_U237_clk),
    .out(_U237_out)
);
assign _U238_in = _U240_out;
_U238_pt__U239 _U238 (
    .in(_U238_in),
    .out(_U238_out)
);
assign _U240_in = 16'(_U228_out + _U331_out);
assign _U240_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U240 (
    .in(_U240_in),
    .clk(_U240_clk),
    .out(_U240_out)
);
assign _U241_in = _U243_out;
_U241_pt__U242 _U241 (
    .in(_U241_in),
    .out(_U241_out)
);
assign _U243_in = 16'(_U252_out + _U393_out);
assign _U243_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U243 (
    .in(_U243_in),
    .clk(_U243_clk),
    .out(_U243_out)
);
assign _U244_in = _U251_out;
_U244_pt__U245 _U244 (
    .in(_U244_in),
    .out(_U244_out)
);
assign _U246_in = 16'(_U378_out * _U359_out);
assign _U246_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U246 (
    .in(_U246_in),
    .clk(_U246_clk),
    .out(_U246_out)
);
assign _U247_in = _U246_out;
assign _U247_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U247 (
    .in(_U247_in),
    .clk(_U247_clk),
    .out(_U247_out)
);
assign _U248_in = _U247_out;
assign _U248_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U248 (
    .in(_U248_in),
    .clk(_U248_clk),
    .out(_U248_out)
);
assign _U249_in = _U248_out;
assign _U249_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U249 (
    .in(_U249_in),
    .clk(_U249_clk),
    .out(_U249_out)
);
assign _U250_in = _U249_out;
assign _U250_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U250 (
    .in(_U250_in),
    .clk(_U250_clk),
    .out(_U250_out)
);
assign _U251_in = _U250_out;
assign _U251_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U251 (
    .in(_U251_in),
    .clk(_U251_clk),
    .out(_U251_out)
);
assign _U252_in = _U255_out;
_U252_pt__U253 _U252 (
    .in(_U252_in),
    .out(_U252_out)
);
assign _U254_in = 16'(_U317_out * _U268_out);
assign _U254_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U254 (
    .in(_U254_in),
    .clk(_U254_clk),
    .out(_U254_out)
);
assign _U255_in = _U254_out;
assign _U255_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U255 (
    .in(_U255_in),
    .clk(_U255_clk),
    .out(_U255_out)
);
assign _U256_in = _U267_out;
_U256_pt__U257 _U256 (
    .in(_U256_in),
    .out(_U256_out)
);
assign _U258_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U258_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U258 (
    .in(_U258_in),
    .clk(_U258_clk),
    .out(_U258_out)
);
assign _U259_in = _U258_out;
assign _U259_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U259 (
    .in(_U259_in),
    .clk(_U259_clk),
    .out(_U259_out)
);
assign _U260_in = _U259_out;
assign _U260_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U260 (
    .in(_U260_in),
    .clk(_U260_clk),
    .out(_U260_out)
);
assign _U261_in = _U260_out;
assign _U261_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U261 (
    .in(_U261_in),
    .clk(_U261_clk),
    .out(_U261_out)
);
assign _U262_in = _U261_out;
assign _U262_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U262 (
    .in(_U262_in),
    .clk(_U262_clk),
    .out(_U262_out)
);
assign _U263_in = _U262_out;
assign _U263_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U263 (
    .in(_U263_in),
    .clk(_U263_clk),
    .out(_U263_out)
);
assign _U264_in = _U263_out;
assign _U264_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U264 (
    .in(_U264_in),
    .clk(_U264_clk),
    .out(_U264_out)
);
assign _U265_in = _U264_out;
assign _U265_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U265 (
    .in(_U265_in),
    .clk(_U265_clk),
    .out(_U265_out)
);
assign _U266_in = _U265_out;
assign _U266_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U266 (
    .in(_U266_in),
    .clk(_U266_clk),
    .out(_U266_out)
);
assign _U267_in = _U266_out;
assign _U267_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U267 (
    .in(_U267_in),
    .clk(_U267_clk),
    .out(_U267_out)
);
assign _U268_in = _U273_out;
_U268_pt__U269 _U268 (
    .in(_U268_in),
    .out(_U268_out)
);
assign _U270_in = in1_hw_input_global_wrapper_stencil[4];
assign _U270_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U270 (
    .in(_U270_in),
    .clk(_U270_clk),
    .out(_U270_out)
);
assign _U271_in = _U270_out;
assign _U271_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U271 (
    .in(_U271_in),
    .clk(_U271_clk),
    .out(_U271_out)
);
assign _U272_in = _U271_out;
assign _U272_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U272 (
    .in(_U272_in),
    .clk(_U272_clk),
    .out(_U272_out)
);
assign _U273_in = _U272_out;
assign _U273_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U273 (
    .in(_U273_in),
    .clk(_U273_clk),
    .out(_U273_out)
);
assign _U274_in = _U279_out;
_U274_pt__U275 _U274 (
    .in(_U274_in),
    .out(_U274_out)
);
assign _U276_in = 16'(_U244_out + _U241_out);
assign _U276_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U276 (
    .in(_U276_in),
    .clk(_U276_clk),
    .out(_U276_out)
);
assign _U277_in = _U276_out;
assign _U277_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U277 (
    .in(_U277_in),
    .clk(_U277_clk),
    .out(_U277_out)
);
assign _U278_in = _U277_out;
assign _U278_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U278 (
    .in(_U278_in),
    .clk(_U278_clk),
    .out(_U278_out)
);
assign _U279_in = _U278_out;
assign _U279_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U279 (
    .in(_U279_in),
    .clk(_U279_clk),
    .out(_U279_out)
);
assign _U280_in = 16'(_U364_out + _U328_out);
_U280_pt__U281 _U280 (
    .in(_U280_in),
    .out(out_conv_stencil)
);
assign _U282_in = _U291_out;
_U282_pt__U283 _U282 (
    .in(_U282_in),
    .out(_U282_out)
);
assign _U284_in = in2_hw_kernel_global_wrapper_stencil[0];
assign _U284_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U284 (
    .in(_U284_in),
    .clk(_U284_clk),
    .out(_U284_out)
);
assign _U285_in = _U284_out;
assign _U285_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U285 (
    .in(_U285_in),
    .clk(_U285_clk),
    .out(_U285_out)
);
assign _U286_in = _U285_out;
assign _U286_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U286 (
    .in(_U286_in),
    .clk(_U286_clk),
    .out(_U286_out)
);
assign _U287_in = _U286_out;
assign _U287_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U287 (
    .in(_U287_in),
    .clk(_U287_clk),
    .out(_U287_out)
);
assign _U288_in = _U287_out;
assign _U288_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U288 (
    .in(_U288_in),
    .clk(_U288_clk),
    .out(_U288_out)
);
assign _U289_in = _U288_out;
assign _U289_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U289 (
    .in(_U289_in),
    .clk(_U289_clk),
    .out(_U289_out)
);
assign _U290_in = _U289_out;
assign _U290_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U290 (
    .in(_U290_in),
    .clk(_U290_clk),
    .out(_U290_out)
);
assign _U291_in = _U290_out;
assign _U291_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U291 (
    .in(_U291_in),
    .clk(_U291_clk),
    .out(_U291_out)
);
assign _U292_in = _U302_out;
_U292_pt__U293 _U292 (
    .in(_U292_in),
    .out(_U292_out)
);
assign _U294_in = in1_hw_input_global_wrapper_stencil[1];
assign _U294_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U294 (
    .in(_U294_in),
    .clk(_U294_clk),
    .out(_U294_out)
);
assign _U295_in = _U294_out;
assign _U295_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U295 (
    .in(_U295_in),
    .clk(_U295_clk),
    .out(_U295_out)
);
assign _U296_in = _U295_out;
assign _U296_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U296 (
    .in(_U296_in),
    .clk(_U296_clk),
    .out(_U296_out)
);
assign _U297_in = _U296_out;
assign _U297_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U297 (
    .in(_U297_in),
    .clk(_U297_clk),
    .out(_U297_out)
);
assign _U298_in = _U297_out;
assign _U298_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U298 (
    .in(_U298_in),
    .clk(_U298_clk),
    .out(_U298_out)
);
assign _U299_in = _U298_out;
assign _U299_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U299 (
    .in(_U299_in),
    .clk(_U299_clk),
    .out(_U299_out)
);
assign _U300_in = _U299_out;
assign _U300_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U300 (
    .in(_U300_in),
    .clk(_U300_clk),
    .out(_U300_out)
);
assign _U301_in = _U300_out;
assign _U301_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U301 (
    .in(_U301_in),
    .clk(_U301_clk),
    .out(_U301_out)
);
assign _U302_in = _U301_out;
assign _U302_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U302 (
    .in(_U302_in),
    .clk(_U302_clk),
    .out(_U302_out)
);
assign _U303_in = _U312_out;
_U303_pt__U304 _U303 (
    .in(_U303_in),
    .out(_U303_out)
);
assign _U305_in = in1_hw_input_global_wrapper_stencil[0];
assign _U305_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U305 (
    .in(_U305_in),
    .clk(_U305_clk),
    .out(_U305_out)
);
assign _U306_in = _U305_out;
assign _U306_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U306 (
    .in(_U306_in),
    .clk(_U306_clk),
    .out(_U306_out)
);
assign _U307_in = _U306_out;
assign _U307_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U307 (
    .in(_U307_in),
    .clk(_U307_clk),
    .out(_U307_out)
);
assign _U308_in = _U307_out;
assign _U308_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U308 (
    .in(_U308_in),
    .clk(_U308_clk),
    .out(_U308_out)
);
assign _U309_in = _U308_out;
assign _U309_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U309 (
    .in(_U309_in),
    .clk(_U309_clk),
    .out(_U309_out)
);
assign _U310_in = _U309_out;
assign _U310_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U310 (
    .in(_U310_in),
    .clk(_U310_clk),
    .out(_U310_out)
);
assign _U311_in = _U310_out;
assign _U311_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U311 (
    .in(_U311_in),
    .clk(_U311_clk),
    .out(_U311_out)
);
assign _U312_in = _U311_out;
assign _U312_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U312 (
    .in(_U312_in),
    .clk(_U312_clk),
    .out(_U312_out)
);
assign _U313_in = _U316_out;
_U313_pt__U314 _U313 (
    .in(_U313_in),
    .out(_U313_out)
);
assign _U315_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U315_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U315 (
    .in(_U315_in),
    .clk(_U315_clk),
    .out(_U315_out)
);
assign _U316_in = _U315_out;
assign _U316_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U316 (
    .in(_U316_in),
    .clk(_U316_clk),
    .out(_U316_out)
);
assign _U317_in = _U322_out;
_U317_pt__U318 _U317 (
    .in(_U317_in),
    .out(_U317_out)
);
assign _U319_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U319_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U319 (
    .in(_U319_in),
    .clk(_U319_clk),
    .out(_U319_out)
);
assign _U320_in = _U319_out;
assign _U320_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U320 (
    .in(_U320_in),
    .clk(_U320_clk),
    .out(_U320_out)
);
assign _U321_in = _U320_out;
assign _U321_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U321 (
    .in(_U321_in),
    .clk(_U321_clk),
    .out(_U321_out)
);
assign _U322_in = _U321_out;
assign _U322_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U322 (
    .in(_U322_in),
    .clk(_U322_clk),
    .out(_U322_out)
);
assign _U323_in = _U327_out;
_U323_pt__U324 _U323 (
    .in(_U323_in),
    .out(_U323_out)
);
assign _U325_in = 16'(_U337_out * _U292_out);
assign _U325_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U325 (
    .in(_U325_in),
    .clk(_U325_clk),
    .out(_U325_out)
);
assign _U326_in = _U325_out;
assign _U326_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U326 (
    .in(_U326_in),
    .clk(_U326_clk),
    .out(_U326_out)
);
assign _U327_in = _U326_out;
assign _U327_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U327 (
    .in(_U327_in),
    .clk(_U327_clk),
    .out(_U327_out)
);
assign _U328_in = _U330_out;
_U328_pt__U329 _U328 (
    .in(_U328_in),
    .out(_U328_out)
);
assign _U330_in = 16'(_U396_out + _U238_out);
assign _U330_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U330 (
    .in(_U330_in),
    .clk(_U330_clk),
    .out(_U330_out)
);
assign _U331_in = _U333_out;
_U331_pt__U332 _U331 (
    .in(_U331_in),
    .out(_U331_out)
);
assign _U333_in = 16'(_U323_out + _U334_out);
assign _U333_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U333 (
    .in(_U333_in),
    .clk(_U333_clk),
    .out(_U333_out)
);
assign _U334_in = _U336_out;
_U334_pt__U335 _U334 (
    .in(_U334_in),
    .out(_U334_out)
);
assign _U336_in = 16'(_U235_out + _U274_out);
assign _U336_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U336 (
    .in(_U336_in),
    .clk(_U336_clk),
    .out(_U336_out)
);
assign _U337_in = _U347_out;
_U337_pt__U338 _U337 (
    .in(_U337_in),
    .out(_U337_out)
);
assign _U339_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U339_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U339 (
    .in(_U339_in),
    .clk(_U339_clk),
    .out(_U339_out)
);
assign _U340_in = _U339_out;
assign _U340_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U340 (
    .in(_U340_in),
    .clk(_U340_clk),
    .out(_U340_out)
);
assign _U341_in = _U340_out;
assign _U341_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U341 (
    .in(_U341_in),
    .clk(_U341_clk),
    .out(_U341_out)
);
assign _U342_in = _U341_out;
assign _U342_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U342 (
    .in(_U342_in),
    .clk(_U342_clk),
    .out(_U342_out)
);
assign _U343_in = _U342_out;
assign _U343_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U343 (
    .in(_U343_in),
    .clk(_U343_clk),
    .out(_U343_out)
);
assign _U344_in = _U343_out;
assign _U344_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U344 (
    .in(_U344_in),
    .clk(_U344_clk),
    .out(_U344_out)
);
assign _U345_in = _U344_out;
assign _U345_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U345 (
    .in(_U345_in),
    .clk(_U345_clk),
    .out(_U345_out)
);
assign _U346_in = _U345_out;
assign _U346_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U346 (
    .in(_U346_in),
    .clk(_U346_clk),
    .out(_U346_out)
);
assign _U347_in = _U346_out;
assign _U347_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U347 (
    .in(_U347_in),
    .clk(_U347_clk),
    .out(_U347_out)
);
assign _U348_in = _U352_out;
_U348_pt__U349 _U348 (
    .in(_U348_in),
    .out(_U348_out)
);
assign _U350_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U350_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U350 (
    .in(_U350_in),
    .clk(_U350_clk),
    .out(_U350_out)
);
assign _U351_in = _U350_out;
assign _U351_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U351 (
    .in(_U351_in),
    .clk(_U351_clk),
    .out(_U351_out)
);
assign _U352_in = _U351_out;
assign _U352_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U352 (
    .in(_U352_in),
    .clk(_U352_clk),
    .out(_U352_out)
);
assign _U353_in = _U356_out;
_U353_pt__U354 _U353 (
    .in(_U353_in),
    .out(_U353_out)
);
assign _U355_in = in1_hw_input_global_wrapper_stencil[5];
assign _U355_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U355 (
    .in(_U355_in),
    .clk(_U355_clk),
    .out(_U355_out)
);
assign _U356_in = _U355_out;
assign _U356_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U356 (
    .in(_U356_in),
    .clk(_U356_clk),
    .out(_U356_out)
);
assign _U357_in = in2_hw_kernel_global_wrapper_stencil[6];
_U357_pt__U358 _U357 (
    .in(_U357_in),
    .out(_U357_out)
);
assign _U359_in = _U361_out;
_U359_pt__U360 _U359 (
    .in(_U359_in),
    .out(_U359_out)
);
assign _U361_in = in1_hw_input_global_wrapper_stencil[3];
assign _U361_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U361 (
    .in(_U361_in),
    .clk(_U361_clk),
    .out(_U361_out)
);
assign _U362_in = in1_hw_input_global_wrapper_stencil[6];
_U362_pt__U363 _U362 (
    .in(_U362_in),
    .out(_U362_out)
);
assign _U364_in = _U377_out;
_U364_pt__U365 _U364 (
    .in(_U364_in),
    .out(_U364_out)
);
assign _U366_in = 16'(_U348_out * _U223_out);
assign _U366_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U366 (
    .in(_U366_in),
    .clk(_U366_clk),
    .out(_U366_out)
);
assign _U367_in = _U366_out;
assign _U367_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U367 (
    .in(_U367_in),
    .clk(_U367_clk),
    .out(_U367_out)
);
assign _U368_in = _U367_out;
assign _U368_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U368 (
    .in(_U368_in),
    .clk(_U368_clk),
    .out(_U368_out)
);
assign _U369_in = _U368_out;
assign _U369_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U369 (
    .in(_U369_in),
    .clk(_U369_clk),
    .out(_U369_out)
);
assign _U370_in = _U369_out;
assign _U370_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U370 (
    .in(_U370_in),
    .clk(_U370_clk),
    .out(_U370_out)
);
assign _U371_in = _U370_out;
assign _U371_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U371 (
    .in(_U371_in),
    .clk(_U371_clk),
    .out(_U371_out)
);
assign _U372_in = _U371_out;
assign _U372_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U372 (
    .in(_U372_in),
    .clk(_U372_clk),
    .out(_U372_out)
);
assign _U373_in = _U372_out;
assign _U373_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U373 (
    .in(_U373_in),
    .clk(_U373_clk),
    .out(_U373_out)
);
assign _U374_in = _U373_out;
assign _U374_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U374 (
    .in(_U374_in),
    .clk(_U374_clk),
    .out(_U374_out)
);
assign _U375_in = _U374_out;
assign _U375_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U375 (
    .in(_U375_in),
    .clk(_U375_clk),
    .out(_U375_out)
);
assign _U376_in = _U375_out;
assign _U376_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U376 (
    .in(_U376_in),
    .clk(_U376_clk),
    .out(_U376_out)
);
assign _U377_in = _U376_out;
assign _U377_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U377 (
    .in(_U377_in),
    .clk(_U377_clk),
    .out(_U377_out)
);
assign _U378_in = _U380_out;
_U378_pt__U379 _U378 (
    .in(_U378_in),
    .out(_U378_out)
);
assign _U380_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U380_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U380 (
    .in(_U380_in),
    .clk(_U380_clk),
    .out(_U380_out)
);
assign _U381_in = _U387_out;
_U381_pt__U382 _U381 (
    .in(_U381_in),
    .out(_U381_out)
);
assign _U383_in = 16'(_U357_out * _U362_out);
assign _U383_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U383 (
    .in(_U383_in),
    .clk(_U383_clk),
    .out(_U383_out)
);
assign _U384_in = _U383_out;
assign _U384_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U384 (
    .in(_U384_in),
    .clk(_U384_clk),
    .out(_U384_out)
);
assign _U385_in = _U384_out;
assign _U385_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U385 (
    .in(_U385_in),
    .clk(_U385_clk),
    .out(_U385_out)
);
assign _U386_in = _U385_out;
assign _U386_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U386 (
    .in(_U386_in),
    .clk(_U386_clk),
    .out(_U386_out)
);
assign _U387_in = _U386_out;
assign _U387_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U387 (
    .in(_U387_in),
    .clk(_U387_clk),
    .out(_U387_out)
);
assign _U388_in = _U392_out;
_U388_pt__U389 _U388 (
    .in(_U388_in),
    .out(_U388_out)
);
assign _U390_in = 16'(_U313_out * _U353_out);
assign _U390_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U390 (
    .in(_U390_in),
    .clk(_U390_clk),
    .out(_U390_out)
);
assign _U391_in = _U390_out;
assign _U391_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U391 (
    .in(_U391_in),
    .clk(_U391_clk),
    .out(_U391_out)
);
assign _U392_in = _U391_out;
assign _U392_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U392 (
    .in(_U392_in),
    .clk(_U392_clk),
    .out(_U392_out)
);
assign _U393_in = _U395_out;
_U393_pt__U394 _U393 (
    .in(_U393_in),
    .out(_U393_out)
);
assign _U395_in = 16'(_U388_out + _U381_out);
assign _U395_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U395 (
    .in(_U395_in),
    .clk(_U395_clk),
    .out(_U395_out)
);
assign _U396_in = _U411_out;
_U396_pt__U397 _U396 (
    .in(_U396_in),
    .out(_U396_out)
);
assign _U398_in = in0_conv_stencil[0];
assign _U398_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U398 (
    .in(_U398_in),
    .clk(_U398_clk),
    .out(_U398_out)
);
assign _U399_in = _U398_out;
assign _U399_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U399 (
    .in(_U399_in),
    .clk(_U399_clk),
    .out(_U399_out)
);
assign _U400_in = _U399_out;
assign _U400_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U400 (
    .in(_U400_in),
    .clk(_U400_clk),
    .out(_U400_out)
);
assign _U401_in = _U400_out;
assign _U401_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U401 (
    .in(_U401_in),
    .clk(_U401_clk),
    .out(_U401_out)
);
assign _U402_in = _U401_out;
assign _U402_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U402 (
    .in(_U402_in),
    .clk(_U402_clk),
    .out(_U402_out)
);
assign _U403_in = _U402_out;
assign _U403_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U403 (
    .in(_U403_in),
    .clk(_U403_clk),
    .out(_U403_out)
);
assign _U404_in = _U403_out;
assign _U404_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U404 (
    .in(_U404_in),
    .clk(_U404_clk),
    .out(_U404_out)
);
assign _U405_in = _U404_out;
assign _U405_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U405 (
    .in(_U405_in),
    .clk(_U405_clk),
    .out(_U405_out)
);
assign _U406_in = _U405_out;
assign _U406_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U406 (
    .in(_U406_in),
    .clk(_U406_clk),
    .out(_U406_out)
);
assign _U407_in = _U406_out;
assign _U407_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U407 (
    .in(_U407_in),
    .clk(_U407_clk),
    .out(_U407_out)
);
assign _U408_in = _U407_out;
assign _U408_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U408 (
    .in(_U408_in),
    .clk(_U408_clk),
    .out(_U408_out)
);
assign _U409_in = _U408_out;
assign _U409_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U409 (
    .in(_U409_in),
    .clk(_U409_clk),
    .out(_U409_out)
);
assign _U410_in = _U409_out;
assign _U410_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U410 (
    .in(_U410_in),
    .clk(_U410_clk),
    .out(_U410_out)
);
assign _U411_in = _U410_out;
assign _U411_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U411 (
    .in(_U411_in),
    .clk(_U411_clk),
    .out(_U411_out)
);
endmodule

module cu_op_hcompute_conv_stencil_4 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
hcompute_conv_stencil_4_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U209_pt__U210 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_hw_kernel_global_wrapper_stencil_pipelined (
    output [15:0] out_hw_kernel_global_wrapper_stencil,
    input [15:0] in0_hw_kernel_stencil [0:0]
);
wire [15:0] _U209_in;
assign _U209_in = in0_hw_kernel_stencil[0];
_U209_pt__U210 _U209 (
    .in(_U209_in),
    .out(out_hw_kernel_global_wrapper_stencil)
);
endmodule

module cu_op_hcompute_hw_kernel_global_wrapper_stencil (
    input clk,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0]
);
wire [15:0] inner_compute_out_hw_kernel_global_wrapper_stencil;
wire [15:0] inner_compute_in0_hw_kernel_stencil [0:0];
assign inner_compute_in0_hw_kernel_stencil[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
hcompute_hw_kernel_global_wrapper_stencil_pipelined inner_compute (
    .out_hw_kernel_global_wrapper_stencil(inner_compute_out_hw_kernel_global_wrapper_stencil),
    .in0_hw_kernel_stencil(inner_compute_in0_hw_kernel_stencil)
);
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = inner_compute_out_hw_kernel_global_wrapper_stencil;
endmodule

module _U206_pt__U207 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U202_pt__U203 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U199_pt__U200 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U182_pt__U183 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U172_pt__U173 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U168_pt__U169 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U164_pt__U165 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U161_pt__U162 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U155_pt__U156 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U148_pt__U149 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U141_pt__U142 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U138_pt__U139 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U133_pt__U134 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U130_pt__U131 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U124_pt__U125 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U11_pt__U12 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U118_pt__U119 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U113_pt__U114 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module _U108_pt__U109 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_5_pipelined (
    input clk,
    input [15:0] in0_conv_stencil [0:0],
    input [15:0] in1_hw_input_global_wrapper_stencil [7:0],
    input [15:0] in2_hw_kernel_global_wrapper_stencil [7:0],
    output [15:0] out_conv_stencil
);
wire [15:0] _U10_in;
wire _U10_clk;
wire [15:0] _U10_out;
wire [15:0] _U100_in;
wire _U100_clk;
wire [15:0] _U100_out;
wire [15:0] _U101_in;
wire _U101_clk;
wire [15:0] _U101_out;
wire [15:0] _U102_in;
wire _U102_clk;
wire [15:0] _U102_out;
wire [15:0] _U103_in;
wire _U103_clk;
wire [15:0] _U103_out;
wire [15:0] _U104_in;
wire _U104_clk;
wire [15:0] _U104_out;
wire [15:0] _U105_in;
wire _U105_clk;
wire [15:0] _U105_out;
wire [15:0] _U106_in;
wire _U106_clk;
wire [15:0] _U106_out;
wire [15:0] _U107_in;
wire _U107_clk;
wire [15:0] _U107_out;
wire [15:0] _U108_in;
wire [15:0] _U108_out;
wire [15:0] _U11_in;
wire [15:0] _U11_out;
wire [15:0] _U110_in;
wire _U110_clk;
wire [15:0] _U110_out;
wire [15:0] _U111_in;
wire _U111_clk;
wire [15:0] _U111_out;
wire [15:0] _U112_in;
wire _U112_clk;
wire [15:0] _U112_out;
wire [15:0] _U113_in;
wire [15:0] _U113_out;
wire [15:0] _U115_in;
wire _U115_clk;
wire [15:0] _U115_out;
wire [15:0] _U116_in;
wire _U116_clk;
wire [15:0] _U116_out;
wire [15:0] _U117_in;
wire _U117_clk;
wire [15:0] _U117_out;
wire [15:0] _U118_in;
wire [15:0] _U118_out;
wire [15:0] _U120_in;
wire _U120_clk;
wire [15:0] _U120_out;
wire [15:0] _U121_in;
wire _U121_clk;
wire [15:0] _U121_out;
wire [15:0] _U122_in;
wire _U122_clk;
wire [15:0] _U122_out;
wire [15:0] _U123_in;
wire _U123_clk;
wire [15:0] _U123_out;
wire [15:0] _U124_in;
wire [15:0] _U124_out;
wire [15:0] _U126_in;
wire _U126_clk;
wire [15:0] _U126_out;
wire [15:0] _U127_in;
wire _U127_clk;
wire [15:0] _U127_out;
wire [15:0] _U128_in;
wire _U128_clk;
wire [15:0] _U128_out;
wire [15:0] _U129_in;
wire _U129_clk;
wire [15:0] _U129_out;
wire [15:0] _U13_in;
wire _U13_clk;
wire [15:0] _U13_out;
wire [15:0] _U130_in;
wire [15:0] _U130_out;
wire [15:0] _U132_in;
wire _U132_clk;
wire [15:0] _U132_out;
wire [15:0] _U133_in;
wire [15:0] _U133_out;
wire [15:0] _U135_in;
wire _U135_clk;
wire [15:0] _U135_out;
wire [15:0] _U136_in;
wire _U136_clk;
wire [15:0] _U136_out;
wire [15:0] _U137_in;
wire _U137_clk;
wire [15:0] _U137_out;
wire [15:0] _U138_in;
wire [15:0] _U138_out;
wire [15:0] _U14_in;
wire _U14_clk;
wire [15:0] _U14_out;
wire [15:0] _U140_in;
wire _U140_clk;
wire [15:0] _U140_out;
wire [15:0] _U141_in;
wire [15:0] _U141_out;
wire [15:0] _U143_in;
wire _U143_clk;
wire [15:0] _U143_out;
wire [15:0] _U144_in;
wire _U144_clk;
wire [15:0] _U144_out;
wire [15:0] _U145_in;
wire _U145_clk;
wire [15:0] _U145_out;
wire [15:0] _U146_in;
wire _U146_clk;
wire [15:0] _U146_out;
wire [15:0] _U147_in;
wire _U147_clk;
wire [15:0] _U147_out;
wire [15:0] _U148_in;
wire [15:0] _U148_out;
wire [15:0] _U15_in;
wire _U15_clk;
wire [15:0] _U15_out;
wire [15:0] _U150_in;
wire _U150_clk;
wire [15:0] _U150_out;
wire [15:0] _U151_in;
wire _U151_clk;
wire [15:0] _U151_out;
wire [15:0] _U152_in;
wire _U152_clk;
wire [15:0] _U152_out;
wire [15:0] _U153_in;
wire _U153_clk;
wire [15:0] _U153_out;
wire [15:0] _U154_in;
wire _U154_clk;
wire [15:0] _U154_out;
wire [15:0] _U155_in;
wire [15:0] _U155_out;
wire [15:0] _U157_in;
wire _U157_clk;
wire [15:0] _U157_out;
wire [15:0] _U158_in;
wire _U158_clk;
wire [15:0] _U158_out;
wire [15:0] _U159_in;
wire _U159_clk;
wire [15:0] _U159_out;
wire [15:0] _U16_in;
wire _U16_clk;
wire [15:0] _U16_out;
wire [15:0] _U160_in;
wire _U160_clk;
wire [15:0] _U160_out;
wire [15:0] _U161_in;
wire [15:0] _U161_out;
wire [15:0] _U163_in;
wire _U163_clk;
wire [15:0] _U163_out;
wire [15:0] _U164_in;
wire [15:0] _U164_out;
wire [15:0] _U166_in;
wire _U166_clk;
wire [15:0] _U166_out;
wire [15:0] _U167_in;
wire _U167_clk;
wire [15:0] _U167_out;
wire [15:0] _U168_in;
wire [15:0] _U168_out;
wire [15:0] _U17_in;
wire _U17_clk;
wire [15:0] _U17_out;
wire [15:0] _U170_in;
wire _U170_clk;
wire [15:0] _U170_out;
wire [15:0] _U171_in;
wire _U171_clk;
wire [15:0] _U171_out;
wire [15:0] _U172_in;
wire [15:0] _U172_out;
wire [15:0] _U174_in;
wire _U174_clk;
wire [15:0] _U174_out;
wire [15:0] _U175_in;
wire _U175_clk;
wire [15:0] _U175_out;
wire [15:0] _U176_in;
wire _U176_clk;
wire [15:0] _U176_out;
wire [15:0] _U177_in;
wire _U177_clk;
wire [15:0] _U177_out;
wire [15:0] _U178_in;
wire _U178_clk;
wire [15:0] _U178_out;
wire [15:0] _U179_in;
wire _U179_clk;
wire [15:0] _U179_out;
wire [15:0] _U18_in;
wire _U18_clk;
wire [15:0] _U18_out;
wire [15:0] _U180_in;
wire _U180_clk;
wire [15:0] _U180_out;
wire [15:0] _U181_in;
wire _U181_clk;
wire [15:0] _U181_out;
wire [15:0] _U182_in;
wire [15:0] _U182_out;
wire [15:0] _U184_in;
wire _U184_clk;
wire [15:0] _U184_out;
wire [15:0] _U185_in;
wire _U185_clk;
wire [15:0] _U185_out;
wire [15:0] _U186_in;
wire _U186_clk;
wire [15:0] _U186_out;
wire [15:0] _U187_in;
wire _U187_clk;
wire [15:0] _U187_out;
wire [15:0] _U188_in;
wire _U188_clk;
wire [15:0] _U188_out;
wire [15:0] _U189_in;
wire _U189_clk;
wire [15:0] _U189_out;
wire [15:0] _U19_in;
wire _U19_clk;
wire [15:0] _U19_out;
wire [15:0] _U190_in;
wire _U190_clk;
wire [15:0] _U190_out;
wire [15:0] _U191_in;
wire _U191_clk;
wire [15:0] _U191_out;
wire [15:0] _U192_in;
wire _U192_clk;
wire [15:0] _U192_out;
wire [15:0] _U193_in;
wire _U193_clk;
wire [15:0] _U193_out;
wire [15:0] _U194_in;
wire _U194_clk;
wire [15:0] _U194_out;
wire [15:0] _U195_in;
wire _U195_clk;
wire [15:0] _U195_out;
wire [15:0] _U196_in;
wire _U196_clk;
wire [15:0] _U196_out;
wire [15:0] _U197_in;
wire _U197_clk;
wire [15:0] _U197_out;
wire [15:0] _U198_in;
wire _U198_clk;
wire [15:0] _U198_out;
wire [15:0] _U199_in;
wire [15:0] _U199_out;
wire [15:0] _U20_in;
wire _U20_clk;
wire [15:0] _U20_out;
wire [15:0] _U201_in;
wire _U201_clk;
wire [15:0] _U201_out;
wire [15:0] _U202_in;
wire [15:0] _U202_out;
wire [15:0] _U204_in;
wire _U204_clk;
wire [15:0] _U204_out;
wire [15:0] _U205_in;
wire _U205_clk;
wire [15:0] _U205_out;
wire [15:0] _U206_in;
wire [15:0] _U206_out;
wire [15:0] _U208_in;
wire _U208_clk;
wire [15:0] _U208_out;
wire [15:0] _U21_in;
wire _U21_clk;
wire [15:0] _U21_out;
wire [15:0] _U22_in;
wire _U22_clk;
wire [15:0] _U22_out;
wire [15:0] _U23_in;
wire _U23_clk;
wire [15:0] _U23_out;
wire [15:0] _U24_in;
wire _U24_clk;
wire [15:0] _U24_out;
wire [15:0] _U25_in;
wire _U25_clk;
wire [15:0] _U25_out;
wire [15:0] _U26_in;
wire _U26_clk;
wire [15:0] _U26_out;
wire [15:0] _U27_in;
wire [15:0] _U27_out;
wire [15:0] _U29_in;
wire _U29_clk;
wire [15:0] _U29_out;
wire [15:0] _U30_in;
wire _U30_clk;
wire [15:0] _U30_out;
wire [15:0] _U31_in;
wire _U31_clk;
wire [15:0] _U31_out;
wire [15:0] _U32_in;
wire _U32_clk;
wire [15:0] _U32_out;
wire [15:0] _U33_in;
wire _U33_clk;
wire [15:0] _U33_out;
wire [15:0] _U34_in;
wire _U34_clk;
wire [15:0] _U34_out;
wire [15:0] _U35_in;
wire _U35_clk;
wire [15:0] _U35_out;
wire [15:0] _U36_in;
wire _U36_clk;
wire [15:0] _U36_out;
wire [15:0] _U37_in;
wire _U37_clk;
wire [15:0] _U37_out;
wire [15:0] _U38_in;
wire _U38_clk;
wire [15:0] _U38_out;
wire [15:0] _U39_in;
wire _U39_clk;
wire [15:0] _U39_out;
wire [15:0] _U40_in;
wire _U40_clk;
wire [15:0] _U40_out;
wire [15:0] _U41_in;
wire [15:0] _U41_out;
wire [15:0] _U43_in;
wire _U43_clk;
wire [15:0] _U43_out;
wire [15:0] _U44_in;
wire [15:0] _U44_out;
wire [15:0] _U46_in;
wire _U46_clk;
wire [15:0] _U46_out;
wire [15:0] _U47_in;
wire [15:0] _U47_out;
wire [15:0] _U49_in;
wire _U49_clk;
wire [15:0] _U49_out;
wire [15:0] _U50_in;
wire _U50_clk;
wire [15:0] _U50_out;
wire [15:0] _U51_in;
wire _U51_clk;
wire [15:0] _U51_out;
wire [15:0] _U52_in;
wire [15:0] _U52_out;
wire [15:0] _U54_in;
wire _U54_clk;
wire [15:0] _U54_out;
wire [15:0] _U55_in;
wire _U55_clk;
wire [15:0] _U55_out;
wire [15:0] _U56_in;
wire _U56_clk;
wire [15:0] _U56_out;
wire [15:0] _U57_in;
wire _U57_clk;
wire [15:0] _U57_out;
wire [15:0] _U58_in;
wire _U58_clk;
wire [15:0] _U58_out;
wire [15:0] _U59_in;
wire _U59_clk;
wire [15:0] _U59_out;
wire [15:0] _U60_in;
wire _U60_clk;
wire [15:0] _U60_out;
wire [15:0] _U61_in;
wire _U61_clk;
wire [15:0] _U61_out;
wire [15:0] _U62_in;
wire _U62_clk;
wire [15:0] _U62_out;
wire [15:0] _U63_in;
wire _U63_clk;
wire [15:0] _U63_out;
wire [15:0] _U64_in;
wire [15:0] _U64_out;
wire [15:0] _U66_in;
wire _U66_clk;
wire [15:0] _U66_out;
wire [15:0] _U67_in;
wire [15:0] _U69_in;
wire [15:0] _U69_out;
wire [15:0] _U71_in;
wire [15:0] _U71_out;
wire [15:0] _U73_in;
wire [15:0] _U73_out;
wire [15:0] _U75_in;
wire _U75_clk;
wire [15:0] _U75_out;
wire [15:0] _U76_in;
wire [15:0] _U76_out;
wire [15:0] _U78_in;
wire _U78_clk;
wire [15:0] _U78_out;
wire [15:0] _U79_in;
wire _U79_clk;
wire [15:0] _U79_out;
wire [15:0] _U8_in;
wire [15:0] _U8_out;
wire [15:0] _U80_in;
wire _U80_clk;
wire [15:0] _U80_out;
wire [15:0] _U81_in;
wire _U81_clk;
wire [15:0] _U81_out;
wire [15:0] _U82_in;
wire _U82_clk;
wire [15:0] _U82_out;
wire [15:0] _U83_in;
wire _U83_clk;
wire [15:0] _U83_out;
wire [15:0] _U84_in;
wire _U84_clk;
wire [15:0] _U84_out;
wire [15:0] _U85_in;
wire _U85_clk;
wire [15:0] _U85_out;
wire [15:0] _U86_in;
wire [15:0] _U86_out;
wire [15:0] _U88_in;
wire _U88_clk;
wire [15:0] _U88_out;
wire [15:0] _U89_in;
wire _U89_clk;
wire [15:0] _U89_out;
wire [15:0] _U90_in;
wire _U90_clk;
wire [15:0] _U90_out;
wire [15:0] _U91_in;
wire _U91_clk;
wire [15:0] _U91_out;
wire [15:0] _U92_in;
wire _U92_clk;
wire [15:0] _U92_out;
wire [15:0] _U93_in;
wire _U93_clk;
wire [15:0] _U93_out;
wire [15:0] _U94_in;
wire _U94_clk;
wire [15:0] _U94_out;
wire [15:0] _U95_in;
wire _U95_clk;
wire [15:0] _U95_out;
wire [15:0] _U96_in;
wire _U96_clk;
wire [15:0] _U96_out;
wire [15:0] _U97_in;
wire [15:0] _U97_out;
wire [15:0] _U99_in;
wire _U99_clk;
wire [15:0] _U99_out;
assign _U10_in = 16'(_U141_out * _U148_out);
assign _U10_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U10 (
    .in(_U10_in),
    .clk(_U10_clk),
    .out(_U10_out)
);
assign _U100_in = _U99_out;
assign _U100_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U100 (
    .in(_U100_in),
    .clk(_U100_clk),
    .out(_U100_out)
);
assign _U101_in = _U100_out;
assign _U101_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U101 (
    .in(_U101_in),
    .clk(_U101_clk),
    .out(_U101_out)
);
assign _U102_in = _U101_out;
assign _U102_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U102 (
    .in(_U102_in),
    .clk(_U102_clk),
    .out(_U102_out)
);
assign _U103_in = _U102_out;
assign _U103_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U103 (
    .in(_U103_in),
    .clk(_U103_clk),
    .out(_U103_out)
);
assign _U104_in = _U103_out;
assign _U104_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U104 (
    .in(_U104_in),
    .clk(_U104_clk),
    .out(_U104_out)
);
assign _U105_in = _U104_out;
assign _U105_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U105 (
    .in(_U105_in),
    .clk(_U105_clk),
    .out(_U105_out)
);
assign _U106_in = _U105_out;
assign _U106_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U106 (
    .in(_U106_in),
    .clk(_U106_clk),
    .out(_U106_out)
);
assign _U107_in = _U106_out;
assign _U107_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U107 (
    .in(_U107_in),
    .clk(_U107_clk),
    .out(_U107_out)
);
assign _U108_in = _U112_out;
_U108_pt__U109 _U108 (
    .in(_U108_in),
    .out(_U108_out)
);
assign _U11_in = _U26_out;
_U11_pt__U12 _U11 (
    .in(_U11_in),
    .out(_U11_out)
);
assign _U110_in = in2_hw_kernel_global_wrapper_stencil[5];
assign _U110_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U110 (
    .in(_U110_in),
    .clk(_U110_clk),
    .out(_U110_out)
);
assign _U111_in = _U110_out;
assign _U111_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U111 (
    .in(_U111_in),
    .clk(_U111_clk),
    .out(_U111_out)
);
assign _U112_in = _U111_out;
assign _U112_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U112 (
    .in(_U112_in),
    .clk(_U112_clk),
    .out(_U112_out)
);
assign _U113_in = _U117_out;
_U113_pt__U114 _U113 (
    .in(_U113_in),
    .out(_U113_out)
);
assign _U115_in = in1_hw_input_global_wrapper_stencil[5];
assign _U115_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U115 (
    .in(_U115_in),
    .clk(_U115_clk),
    .out(_U115_out)
);
assign _U116_in = _U115_out;
assign _U116_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U116 (
    .in(_U116_in),
    .clk(_U116_clk),
    .out(_U116_out)
);
assign _U117_in = _U116_out;
assign _U117_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U117 (
    .in(_U117_in),
    .clk(_U117_clk),
    .out(_U117_out)
);
assign _U118_in = _U123_out;
_U118_pt__U119 _U118 (
    .in(_U118_in),
    .out(_U118_out)
);
assign _U120_in = in2_hw_kernel_global_wrapper_stencil[6];
assign _U120_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U120 (
    .in(_U120_in),
    .clk(_U120_clk),
    .out(_U120_out)
);
assign _U121_in = _U120_out;
assign _U121_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U121 (
    .in(_U121_in),
    .clk(_U121_clk),
    .out(_U121_out)
);
assign _U122_in = _U121_out;
assign _U122_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U122 (
    .in(_U122_in),
    .clk(_U122_clk),
    .out(_U122_out)
);
assign _U123_in = _U122_out;
assign _U123_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U123 (
    .in(_U123_in),
    .clk(_U123_clk),
    .out(_U123_out)
);
assign _U124_in = _U129_out;
_U124_pt__U125 _U124 (
    .in(_U124_in),
    .out(_U124_out)
);
assign _U126_in = in1_hw_input_global_wrapper_stencil[6];
assign _U126_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U126 (
    .in(_U126_in),
    .clk(_U126_clk),
    .out(_U126_out)
);
assign _U127_in = _U126_out;
assign _U127_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U127 (
    .in(_U127_in),
    .clk(_U127_clk),
    .out(_U127_out)
);
assign _U128_in = _U127_out;
assign _U128_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U128 (
    .in(_U128_in),
    .clk(_U128_clk),
    .out(_U128_out)
);
assign _U129_in = _U128_out;
assign _U129_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U129 (
    .in(_U129_in),
    .clk(_U129_clk),
    .out(_U129_out)
);
assign _U13_in = in0_conv_stencil[0];
assign _U13_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U13 (
    .in(_U13_in),
    .clk(_U13_clk),
    .out(_U13_out)
);
assign _U130_in = _U132_out;
_U130_pt__U131 _U130 (
    .in(_U130_in),
    .out(_U130_out)
);
assign _U132_in = 16'(_U52_out + _U64_out);
assign _U132_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U132 (
    .in(_U132_in),
    .clk(_U132_clk),
    .out(_U132_out)
);
assign _U133_in = _U137_out;
_U133_pt__U134 _U133 (
    .in(_U133_in),
    .out(_U133_out)
);
assign _U135_in = 16'(_U172_out * _U76_out);
assign _U135_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U135 (
    .in(_U135_in),
    .clk(_U135_clk),
    .out(_U135_out)
);
assign _U136_in = _U135_out;
assign _U136_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U136 (
    .in(_U136_in),
    .clk(_U136_clk),
    .out(_U136_out)
);
assign _U137_in = _U136_out;
assign _U137_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U137 (
    .in(_U137_in),
    .clk(_U137_clk),
    .out(_U137_out)
);
assign _U138_in = _U140_out;
_U138_pt__U139 _U138 (
    .in(_U138_in),
    .out(_U138_out)
);
assign _U14_in = _U13_out;
assign _U14_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U14 (
    .in(_U14_in),
    .clk(_U14_clk),
    .out(_U14_out)
);
assign _U140_in = 16'(_U44_out + _U47_out);
assign _U140_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U140 (
    .in(_U140_in),
    .clk(_U140_clk),
    .out(_U140_out)
);
assign _U141_in = _U147_out;
_U141_pt__U142 _U141 (
    .in(_U141_in),
    .out(_U141_out)
);
assign _U143_in = in2_hw_kernel_global_wrapper_stencil[7];
assign _U143_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U143 (
    .in(_U143_in),
    .clk(_U143_clk),
    .out(_U143_out)
);
assign _U144_in = _U143_out;
assign _U144_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U144 (
    .in(_U144_in),
    .clk(_U144_clk),
    .out(_U144_out)
);
assign _U145_in = _U144_out;
assign _U145_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U145 (
    .in(_U145_in),
    .clk(_U145_clk),
    .out(_U145_out)
);
assign _U146_in = _U145_out;
assign _U146_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U146 (
    .in(_U146_in),
    .clk(_U146_clk),
    .out(_U146_out)
);
assign _U147_in = _U146_out;
assign _U147_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U147 (
    .in(_U147_in),
    .clk(_U147_clk),
    .out(_U147_out)
);
assign _U148_in = _U154_out;
_U148_pt__U149 _U148 (
    .in(_U148_in),
    .out(_U148_out)
);
assign _U15_in = _U14_out;
assign _U15_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U15 (
    .in(_U15_in),
    .clk(_U15_clk),
    .out(_U15_out)
);
assign _U150_in = in1_hw_input_global_wrapper_stencil[7];
assign _U150_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U150 (
    .in(_U150_in),
    .clk(_U150_clk),
    .out(_U150_out)
);
assign _U151_in = _U150_out;
assign _U151_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U151 (
    .in(_U151_in),
    .clk(_U151_clk),
    .out(_U151_out)
);
assign _U152_in = _U151_out;
assign _U152_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U152 (
    .in(_U152_in),
    .clk(_U152_clk),
    .out(_U152_out)
);
assign _U153_in = _U152_out;
assign _U153_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U153 (
    .in(_U153_in),
    .clk(_U153_clk),
    .out(_U153_out)
);
assign _U154_in = _U153_out;
assign _U154_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U154 (
    .in(_U154_in),
    .clk(_U154_clk),
    .out(_U154_out)
);
assign _U155_in = _U160_out;
_U155_pt__U156 _U155 (
    .in(_U155_in),
    .out(_U155_out)
);
assign _U157_in = 16'(_U108_out * _U113_out);
assign _U157_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U157 (
    .in(_U157_in),
    .clk(_U157_clk),
    .out(_U157_out)
);
assign _U158_in = _U157_out;
assign _U158_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U158 (
    .in(_U158_in),
    .clk(_U158_clk),
    .out(_U158_out)
);
assign _U159_in = _U158_out;
assign _U159_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U159 (
    .in(_U159_in),
    .clk(_U159_clk),
    .out(_U159_out)
);
assign _U16_in = _U15_out;
assign _U16_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U16 (
    .in(_U16_in),
    .clk(_U16_clk),
    .out(_U16_out)
);
assign _U160_in = _U159_out;
assign _U160_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U160 (
    .in(_U160_in),
    .clk(_U160_clk),
    .out(_U160_out)
);
assign _U161_in = _U163_out;
_U161_pt__U162 _U161 (
    .in(_U161_in),
    .out(_U161_out)
);
assign _U163_in = in1_hw_input_global_wrapper_stencil[1];
assign _U163_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U163 (
    .in(_U163_in),
    .clk(_U163_clk),
    .out(_U163_out)
);
assign _U164_in = _U167_out;
_U164_pt__U165 _U164 (
    .in(_U164_in),
    .out(_U164_out)
);
assign _U166_in = in2_hw_kernel_global_wrapper_stencil[2];
assign _U166_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U166 (
    .in(_U166_in),
    .clk(_U166_clk),
    .out(_U166_out)
);
assign _U167_in = _U166_out;
assign _U167_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U167 (
    .in(_U167_in),
    .clk(_U167_clk),
    .out(_U167_out)
);
assign _U168_in = _U171_out;
_U168_pt__U169 _U168 (
    .in(_U168_in),
    .out(_U168_out)
);
assign _U17_in = _U16_out;
assign _U17_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U17 (
    .in(_U17_in),
    .clk(_U17_clk),
    .out(_U17_out)
);
assign _U170_in = in1_hw_input_global_wrapper_stencil[2];
assign _U170_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U170 (
    .in(_U170_in),
    .clk(_U170_clk),
    .out(_U170_out)
);
assign _U171_in = _U170_out;
assign _U171_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U171 (
    .in(_U171_in),
    .clk(_U171_clk),
    .out(_U171_out)
);
assign _U172_in = _U181_out;
_U172_pt__U173 _U172 (
    .in(_U172_in),
    .out(_U172_out)
);
assign _U174_in = in2_hw_kernel_global_wrapper_stencil[3];
assign _U174_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U174 (
    .in(_U174_in),
    .clk(_U174_clk),
    .out(_U174_out)
);
assign _U175_in = _U174_out;
assign _U175_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U175 (
    .in(_U175_in),
    .clk(_U175_clk),
    .out(_U175_out)
);
assign _U176_in = _U175_out;
assign _U176_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U176 (
    .in(_U176_in),
    .clk(_U176_clk),
    .out(_U176_out)
);
assign _U177_in = _U176_out;
assign _U177_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U177 (
    .in(_U177_in),
    .clk(_U177_clk),
    .out(_U177_out)
);
assign _U178_in = _U177_out;
assign _U178_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U178 (
    .in(_U178_in),
    .clk(_U178_clk),
    .out(_U178_out)
);
assign _U179_in = _U178_out;
assign _U179_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U179 (
    .in(_U179_in),
    .clk(_U179_clk),
    .out(_U179_out)
);
assign _U18_in = _U17_out;
assign _U18_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U18 (
    .in(_U18_in),
    .clk(_U18_clk),
    .out(_U18_out)
);
assign _U180_in = _U179_out;
assign _U180_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U180 (
    .in(_U180_in),
    .clk(_U180_clk),
    .out(_U180_out)
);
assign _U181_in = _U180_out;
assign _U181_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U181 (
    .in(_U181_in),
    .clk(_U181_clk),
    .out(_U181_out)
);
assign _U182_in = _U198_out;
_U182_pt__U183 _U182 (
    .in(_U182_in),
    .out(_U182_out)
);
assign _U184_in = 16'(_U69_out * _U71_out);
assign _U184_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U184 (
    .in(_U184_in),
    .clk(_U184_clk),
    .out(_U184_out)
);
assign _U185_in = _U184_out;
assign _U185_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U185 (
    .in(_U185_in),
    .clk(_U185_clk),
    .out(_U185_out)
);
assign _U186_in = _U185_out;
assign _U186_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U186 (
    .in(_U186_in),
    .clk(_U186_clk),
    .out(_U186_out)
);
assign _U187_in = _U186_out;
assign _U187_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U187 (
    .in(_U187_in),
    .clk(_U187_clk),
    .out(_U187_out)
);
assign _U188_in = _U187_out;
assign _U188_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U188 (
    .in(_U188_in),
    .clk(_U188_clk),
    .out(_U188_out)
);
assign _U189_in = _U188_out;
assign _U189_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U189 (
    .in(_U189_in),
    .clk(_U189_clk),
    .out(_U189_out)
);
assign _U19_in = _U18_out;
assign _U19_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U19 (
    .in(_U19_in),
    .clk(_U19_clk),
    .out(_U19_out)
);
assign _U190_in = _U189_out;
assign _U190_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U190 (
    .in(_U190_in),
    .clk(_U190_clk),
    .out(_U190_out)
);
assign _U191_in = _U190_out;
assign _U191_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U191 (
    .in(_U191_in),
    .clk(_U191_clk),
    .out(_U191_out)
);
assign _U192_in = _U191_out;
assign _U192_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U192 (
    .in(_U192_in),
    .clk(_U192_clk),
    .out(_U192_out)
);
assign _U193_in = _U192_out;
assign _U193_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U193 (
    .in(_U193_in),
    .clk(_U193_clk),
    .out(_U193_out)
);
assign _U194_in = _U193_out;
assign _U194_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U194 (
    .in(_U194_in),
    .clk(_U194_clk),
    .out(_U194_out)
);
assign _U195_in = _U194_out;
assign _U195_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U195 (
    .in(_U195_in),
    .clk(_U195_clk),
    .out(_U195_out)
);
assign _U196_in = _U195_out;
assign _U196_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U196 (
    .in(_U196_in),
    .clk(_U196_clk),
    .out(_U196_out)
);
assign _U197_in = _U196_out;
assign _U197_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U197 (
    .in(_U197_in),
    .clk(_U197_clk),
    .out(_U197_out)
);
assign _U198_in = _U197_out;
assign _U198_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U198 (
    .in(_U198_in),
    .clk(_U198_clk),
    .out(_U198_out)
);
assign _U199_in = _U201_out;
_U199_pt__U200 _U199 (
    .in(_U199_in),
    .out(_U199_out)
);
assign _U20_in = _U19_out;
assign _U20_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U20 (
    .in(_U20_in),
    .clk(_U20_clk),
    .out(_U20_out)
);
assign _U201_in = 16'(_U11_out + _U41_out);
assign _U201_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U201 (
    .in(_U201_in),
    .clk(_U201_clk),
    .out(_U201_out)
);
assign _U202_in = _U205_out;
_U202_pt__U203 _U202 (
    .in(_U202_in),
    .out(_U202_out)
);
assign _U204_in = 16'(_U118_out * _U124_out);
assign _U204_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U204 (
    .in(_U204_in),
    .clk(_U204_clk),
    .out(_U204_out)
);
assign _U205_in = _U204_out;
assign _U205_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U205 (
    .in(_U205_in),
    .clk(_U205_clk),
    .out(_U205_out)
);
assign _U206_in = _U208_out;
_U206_pt__U207 _U206 (
    .in(_U206_in),
    .out(_U206_out)
);
assign _U208_in = 16'(_U202_out + _U8_out);
assign _U208_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U208 (
    .in(_U208_in),
    .clk(_U208_clk),
    .out(_U208_out)
);
assign _U21_in = _U20_out;
assign _U21_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U21 (
    .in(_U21_in),
    .clk(_U21_clk),
    .out(_U21_out)
);
assign _U22_in = _U21_out;
assign _U22_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U22 (
    .in(_U22_in),
    .clk(_U22_clk),
    .out(_U22_out)
);
assign _U23_in = _U22_out;
assign _U23_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U23 (
    .in(_U23_in),
    .clk(_U23_clk),
    .out(_U23_out)
);
assign _U24_in = _U23_out;
assign _U24_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U24 (
    .in(_U24_in),
    .clk(_U24_clk),
    .out(_U24_out)
);
assign _U25_in = _U24_out;
assign _U25_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U25 (
    .in(_U25_in),
    .clk(_U25_clk),
    .out(_U25_out)
);
assign _U26_in = _U25_out;
assign _U26_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U26 (
    .in(_U26_in),
    .clk(_U26_clk),
    .out(_U26_out)
);
assign _U27_in = _U40_out;
_U27_pt__U28 _U27 (
    .in(_U27_in),
    .out(_U27_out)
);
assign _U29_in = 16'(_U73_out * _U161_out);
assign _U29_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U29 (
    .in(_U29_in),
    .clk(_U29_clk),
    .out(_U29_out)
);
assign _U30_in = _U29_out;
assign _U30_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U30 (
    .in(_U30_in),
    .clk(_U30_clk),
    .out(_U30_out)
);
assign _U31_in = _U30_out;
assign _U31_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U31 (
    .in(_U31_in),
    .clk(_U31_clk),
    .out(_U31_out)
);
assign _U32_in = _U31_out;
assign _U32_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U32 (
    .in(_U32_in),
    .clk(_U32_clk),
    .out(_U32_out)
);
assign _U33_in = _U32_out;
assign _U33_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U33 (
    .in(_U33_in),
    .clk(_U33_clk),
    .out(_U33_out)
);
assign _U34_in = _U33_out;
assign _U34_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U34 (
    .in(_U34_in),
    .clk(_U34_clk),
    .out(_U34_out)
);
assign _U35_in = _U34_out;
assign _U35_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U35 (
    .in(_U35_in),
    .clk(_U35_clk),
    .out(_U35_out)
);
assign _U36_in = _U35_out;
assign _U36_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U36 (
    .in(_U36_in),
    .clk(_U36_clk),
    .out(_U36_out)
);
assign _U37_in = _U36_out;
assign _U37_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U37 (
    .in(_U37_in),
    .clk(_U37_clk),
    .out(_U37_out)
);
assign _U38_in = _U37_out;
assign _U38_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U38 (
    .in(_U38_in),
    .clk(_U38_clk),
    .out(_U38_out)
);
assign _U39_in = _U38_out;
assign _U39_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U39 (
    .in(_U39_in),
    .clk(_U39_clk),
    .out(_U39_out)
);
assign _U40_in = _U39_out;
assign _U40_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U40 (
    .in(_U40_in),
    .clk(_U40_clk),
    .out(_U40_out)
);
assign _U41_in = _U43_out;
_U41_pt__U42 _U41 (
    .in(_U41_in),
    .out(_U41_out)
);
assign _U43_in = 16'(_U27_out + _U130_out);
assign _U43_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U43 (
    .in(_U43_in),
    .clk(_U43_clk),
    .out(_U43_out)
);
assign _U44_in = _U46_out;
_U44_pt__U45 _U44 (
    .in(_U44_in),
    .out(_U44_out)
);
assign _U46_in = 16'(_U86_out * _U97_out);
assign _U46_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U46 (
    .in(_U46_in),
    .clk(_U46_clk),
    .out(_U46_out)
);
assign _U47_in = _U51_out;
_U47_pt__U48 _U47 (
    .in(_U47_in),
    .out(_U47_out)
);
assign _U49_in = 16'(_U155_out + _U206_out);
assign _U49_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U49 (
    .in(_U49_in),
    .clk(_U49_clk),
    .out(_U49_out)
);
assign _U50_in = _U49_out;
assign _U50_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U50 (
    .in(_U50_in),
    .clk(_U50_clk),
    .out(_U50_out)
);
assign _U51_in = _U50_out;
assign _U51_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U51 (
    .in(_U51_in),
    .clk(_U51_clk),
    .out(_U51_out)
);
assign _U52_in = _U63_out;
_U52_pt__U53 _U52 (
    .in(_U52_in),
    .out(_U52_out)
);
assign _U54_in = 16'(_U164_out * _U168_out);
assign _U54_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U54 (
    .in(_U54_in),
    .clk(_U54_clk),
    .out(_U54_out)
);
assign _U55_in = _U54_out;
assign _U55_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U55 (
    .in(_U55_in),
    .clk(_U55_clk),
    .out(_U55_out)
);
assign _U56_in = _U55_out;
assign _U56_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U56 (
    .in(_U56_in),
    .clk(_U56_clk),
    .out(_U56_out)
);
assign _U57_in = _U56_out;
assign _U57_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U57 (
    .in(_U57_in),
    .clk(_U57_clk),
    .out(_U57_out)
);
assign _U58_in = _U57_out;
assign _U58_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U58 (
    .in(_U58_in),
    .clk(_U58_clk),
    .out(_U58_out)
);
assign _U59_in = _U58_out;
assign _U59_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U59 (
    .in(_U59_in),
    .clk(_U59_clk),
    .out(_U59_out)
);
assign _U60_in = _U59_out;
assign _U60_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U60 (
    .in(_U60_in),
    .clk(_U60_clk),
    .out(_U60_out)
);
assign _U61_in = _U60_out;
assign _U61_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U61 (
    .in(_U61_in),
    .clk(_U61_clk),
    .out(_U61_out)
);
assign _U62_in = _U61_out;
assign _U62_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U62 (
    .in(_U62_in),
    .clk(_U62_clk),
    .out(_U62_out)
);
assign _U63_in = _U62_out;
assign _U63_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U63 (
    .in(_U63_in),
    .clk(_U63_clk),
    .out(_U63_out)
);
assign _U64_in = _U66_out;
_U64_pt__U65 _U64 (
    .in(_U64_in),
    .out(_U64_out)
);
assign _U66_in = 16'(_U133_out + _U138_out);
assign _U66_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U66 (
    .in(_U66_in),
    .clk(_U66_clk),
    .out(_U66_out)
);
assign _U67_in = 16'(_U182_out + _U199_out);
_U67_pt__U68 _U67 (
    .in(_U67_in),
    .out(out_conv_stencil)
);
assign _U69_in = in2_hw_kernel_global_wrapper_stencil[0];
_U69_pt__U70 _U69 (
    .in(_U69_in),
    .out(_U69_out)
);
assign _U71_in = in1_hw_input_global_wrapper_stencil[0];
_U71_pt__U72 _U71 (
    .in(_U71_in),
    .out(_U71_out)
);
assign _U73_in = _U75_out;
_U73_pt__U74 _U73 (
    .in(_U73_in),
    .out(_U73_out)
);
assign _U75_in = in2_hw_kernel_global_wrapper_stencil[1];
assign _U75_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U75 (
    .in(_U75_in),
    .clk(_U75_clk),
    .out(_U75_out)
);
assign _U76_in = _U85_out;
_U76_pt__U77 _U76 (
    .in(_U76_in),
    .out(_U76_out)
);
assign _U78_in = in1_hw_input_global_wrapper_stencil[3];
assign _U78_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U78 (
    .in(_U78_in),
    .clk(_U78_clk),
    .out(_U78_out)
);
assign _U79_in = _U78_out;
assign _U79_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U79 (
    .in(_U79_in),
    .clk(_U79_clk),
    .out(_U79_out)
);
assign _U8_in = _U10_out;
_U8_pt__U9 _U8 (
    .in(_U8_in),
    .out(_U8_out)
);
assign _U80_in = _U79_out;
assign _U80_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U80 (
    .in(_U80_in),
    .clk(_U80_clk),
    .out(_U80_out)
);
assign _U81_in = _U80_out;
assign _U81_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U81 (
    .in(_U81_in),
    .clk(_U81_clk),
    .out(_U81_out)
);
assign _U82_in = _U81_out;
assign _U82_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U82 (
    .in(_U82_in),
    .clk(_U82_clk),
    .out(_U82_out)
);
assign _U83_in = _U82_out;
assign _U83_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U83 (
    .in(_U83_in),
    .clk(_U83_clk),
    .out(_U83_out)
);
assign _U84_in = _U83_out;
assign _U84_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U84 (
    .in(_U84_in),
    .clk(_U84_clk),
    .out(_U84_out)
);
assign _U85_in = _U84_out;
assign _U85_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U85 (
    .in(_U85_in),
    .clk(_U85_clk),
    .out(_U85_out)
);
assign _U86_in = _U96_out;
_U86_pt__U87 _U86 (
    .in(_U86_in),
    .out(_U86_out)
);
assign _U88_in = in2_hw_kernel_global_wrapper_stencil[4];
assign _U88_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U88 (
    .in(_U88_in),
    .clk(_U88_clk),
    .out(_U88_out)
);
assign _U89_in = _U88_out;
assign _U89_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U89 (
    .in(_U89_in),
    .clk(_U89_clk),
    .out(_U89_out)
);
assign _U90_in = _U89_out;
assign _U90_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U90 (
    .in(_U90_in),
    .clk(_U90_clk),
    .out(_U90_out)
);
assign _U91_in = _U90_out;
assign _U91_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U91 (
    .in(_U91_in),
    .clk(_U91_clk),
    .out(_U91_out)
);
assign _U92_in = _U91_out;
assign _U92_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U92 (
    .in(_U92_in),
    .clk(_U92_clk),
    .out(_U92_out)
);
assign _U93_in = _U92_out;
assign _U93_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U93 (
    .in(_U93_in),
    .clk(_U93_clk),
    .out(_U93_out)
);
assign _U94_in = _U93_out;
assign _U94_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U94 (
    .in(_U94_in),
    .clk(_U94_clk),
    .out(_U94_out)
);
assign _U95_in = _U94_out;
assign _U95_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U95 (
    .in(_U95_in),
    .clk(_U95_clk),
    .out(_U95_out)
);
assign _U96_in = _U95_out;
assign _U96_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U96 (
    .in(_U96_in),
    .clk(_U96_clk),
    .out(_U96_out)
);
assign _U97_in = _U107_out;
_U97_pt__U98 _U97 (
    .in(_U97_in),
    .out(_U97_out)
);
assign _U99_in = in1_hw_input_global_wrapper_stencil[4];
assign _U99_clk = clk;
mantle_reg__has_clrFalse__has_enFalse__has_rstFalse__width16 #(
    .init(16'h0000)
) _U99 (
    .in(_U99_in),
    .clk(_U99_clk),
    .out(_U99_out)
);
endmodule

module cu_op_hcompute_conv_stencil_5 (
    input clk,
    input [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0],
    input [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    input [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0],
    output [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0]
);
wire inner_compute_clk;
wire [15:0] inner_compute_in0_conv_stencil [0:0];
wire [15:0] inner_compute_in1_hw_input_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_in2_hw_kernel_global_wrapper_stencil [7:0];
wire [15:0] inner_compute_out_conv_stencil;
assign inner_compute_clk = clk;
assign inner_compute_in0_conv_stencil[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in1_hw_input_global_wrapper_stencil[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in1_hw_input_global_wrapper_stencil[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in1_hw_input_global_wrapper_stencil[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in1_hw_input_global_wrapper_stencil[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in1_hw_input_global_wrapper_stencil[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in1_hw_input_global_wrapper_stencil[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in1_hw_input_global_wrapper_stencil[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in1_hw_input_global_wrapper_stencil[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign inner_compute_in2_hw_kernel_global_wrapper_stencil[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
hcompute_conv_stencil_5_pipelined inner_compute (
    .clk(inner_compute_clk),
    .in0_conv_stencil(inner_compute_in0_conv_stencil),
    .in1_hw_input_global_wrapper_stencil(inner_compute_in1_hw_input_global_wrapper_stencil),
    .in2_hw_kernel_global_wrapper_stencil(inner_compute_in2_hw_kernel_global_wrapper_stencil),
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = inner_compute_out_conv_stencil;
endmodule

module _U0_pt__U1 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module hcompute_conv_stencil_pipelined (
    output [15:0] out_conv_stencil
);
wire [15:0] _U0_in;
assign _U0_in = 16'h0000;
_U0_pt__U1 _U0 (
    .in(_U0_in),
    .out(out_conv_stencil)
);
endmodule

module cu_op_hcompute_conv_stencil (
    input clk,
    output [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0]
);
wire [15:0] inner_compute_out_conv_stencil;
hcompute_conv_stencil_pipelined inner_compute (
    .out_conv_stencil(inner_compute_out_conv_stencil)
);
assign conv_stencil_op_hcompute_conv_stencil_write[0] = inner_compute_out_conv_stencil;
endmodule

module resnet (
    input clk,
    input rst_n,
    input flush,
    output hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en,
    input [15:0] hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0],
    output hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en,
    input [15:0] hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0],
    output hw_output_stencil_op_hcompute_hw_output_stencil_write_valid,
    output [15:0] hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0]
);
wire arr__U104_clk;
wire [15:0] arr__U104_in [3:0];
wire [15:0] arr__U104_out [3:0];
wire arr__U114_clk;
wire [15:0] arr__U114_in [3:0];
wire [15:0] arr__U114_out [3:0];
wire arr__U120_clk;
wire [15:0] arr__U120_in [3:0];
wire [15:0] arr__U120_out [3:0];
wire arr__U162_clk;
wire [15:0] arr__U162_in [4:0];
wire [15:0] arr__U162_out [4:0];
wire arr__U169_clk;
wire [15:0] arr__U169_in [4:0];
wire [15:0] arr__U169_out [4:0];
wire arr__U195_clk;
wire [15:0] arr__U195_in [4:0];
wire [15:0] arr__U195_out [4:0];
wire arr__U202_clk;
wire [15:0] arr__U202_in [4:0];
wire [15:0] arr__U202_out [4:0];
wire arr__U209_clk;
wire [15:0] arr__U209_in [4:0];
wire [15:0] arr__U209_out [4:0];
wire arr__U216_clk;
wire [15:0] arr__U216_in [4:0];
wire [15:0] arr__U216_out [4:0];
wire arr__U223_clk;
wire [15:0] arr__U223_in [4:0];
wire [15:0] arr__U223_out [4:0];
wire arr__U230_clk;
wire [15:0] arr__U230_in [4:0];
wire [15:0] arr__U230_out [4:0];
wire arr__U237_clk;
wire [15:0] arr__U237_in [4:0];
wire [15:0] arr__U237_out [4:0];
wire arr__U244_clk;
wire [15:0] arr__U244_in [4:0];
wire [15:0] arr__U244_out [4:0];
wire arr__U251_clk;
wire [15:0] arr__U251_in [4:0];
wire [15:0] arr__U251_out [4:0];
wire arr__U258_clk;
wire [15:0] arr__U258_in [4:0];
wire [15:0] arr__U258_out [4:0];
wire arr__U265_clk;
wire [15:0] arr__U265_in [4:0];
wire [15:0] arr__U265_out [4:0];
wire arr__U272_clk;
wire [15:0] arr__U272_in [4:0];
wire [15:0] arr__U272_out [4:0];
wire arr__U279_clk;
wire [15:0] arr__U279_in [4:0];
wire [15:0] arr__U279_out [4:0];
wire arr__U286_clk;
wire [15:0] arr__U286_in [4:0];
wire [15:0] arr__U286_out [4:0];
wire arr__U293_clk;
wire [15:0] arr__U293_in [4:0];
wire [15:0] arr__U293_out [4:0];
wire arr__U300_clk;
wire [15:0] arr__U300_in [4:0];
wire [15:0] arr__U300_out [4:0];
wire arr__U307_clk;
wire [15:0] arr__U307_in [4:0];
wire [15:0] arr__U307_out [4:0];
wire arr__U386_clk;
wire [15:0] arr__U386_in [4:0];
wire [15:0] arr__U386_out [4:0];
wire arr__U393_clk;
wire [15:0] arr__U393_in [4:0];
wire [15:0] arr__U393_out [4:0];
wire arr__U419_clk;
wire [15:0] arr__U419_in [4:0];
wire [15:0] arr__U419_out [4:0];
wire arr__U426_clk;
wire [15:0] arr__U426_in [4:0];
wire [15:0] arr__U426_out [4:0];
wire arr__U433_clk;
wire [15:0] arr__U433_in [4:0];
wire [15:0] arr__U433_out [4:0];
wire arr__U440_clk;
wire [15:0] arr__U440_in [4:0];
wire [15:0] arr__U440_out [4:0];
wire arr__U447_clk;
wire [15:0] arr__U447_in [4:0];
wire [15:0] arr__U447_out [4:0];
wire arr__U454_clk;
wire [15:0] arr__U454_in [4:0];
wire [15:0] arr__U454_out [4:0];
wire arr__U461_clk;
wire [15:0] arr__U461_in [4:0];
wire [15:0] arr__U461_out [4:0];
wire arr__U468_clk;
wire [15:0] arr__U468_in [4:0];
wire [15:0] arr__U468_out [4:0];
wire arr__U475_clk;
wire [15:0] arr__U475_in [4:0];
wire [15:0] arr__U475_out [4:0];
wire arr__U482_clk;
wire [15:0] arr__U482_in [4:0];
wire [15:0] arr__U482_out [4:0];
wire arr__U489_clk;
wire [15:0] arr__U489_in [4:0];
wire [15:0] arr__U489_out [4:0];
wire arr__U496_clk;
wire [15:0] arr__U496_in [4:0];
wire [15:0] arr__U496_out [4:0];
wire arr__U503_clk;
wire [15:0] arr__U503_in [4:0];
wire [15:0] arr__U503_out [4:0];
wire arr__U510_clk;
wire [15:0] arr__U510_in [4:0];
wire [15:0] arr__U510_out [4:0];
wire arr__U517_clk;
wire [15:0] arr__U517_in [4:0];
wire [15:0] arr__U517_out [4:0];
wire arr__U524_clk;
wire [15:0] arr__U524_in [4:0];
wire [15:0] arr__U524_out [4:0];
wire arr__U531_clk;
wire [15:0] arr__U531_in [4:0];
wire [15:0] arr__U531_out [4:0];
wire arr__U574_clk;
wire [15:0] arr__U574_in [4:0];
wire [15:0] arr__U574_out [4:0];
wire arr__U581_clk;
wire [15:0] arr__U581_in [4:0];
wire [15:0] arr__U581_out [4:0];
wire arr__U607_clk;
wire [15:0] arr__U607_in [4:0];
wire [15:0] arr__U607_out [4:0];
wire arr__U614_clk;
wire [15:0] arr__U614_in [4:0];
wire [15:0] arr__U614_out [4:0];
wire arr__U621_clk;
wire [15:0] arr__U621_in [4:0];
wire [15:0] arr__U621_out [4:0];
wire arr__U628_clk;
wire [15:0] arr__U628_in [4:0];
wire [15:0] arr__U628_out [4:0];
wire arr__U635_clk;
wire [15:0] arr__U635_in [4:0];
wire [15:0] arr__U635_out [4:0];
wire arr__U642_clk;
wire [15:0] arr__U642_in [4:0];
wire [15:0] arr__U642_out [4:0];
wire arr__U649_clk;
wire [15:0] arr__U649_in [4:0];
wire [15:0] arr__U649_out [4:0];
wire arr__U656_clk;
wire [15:0] arr__U656_in [4:0];
wire [15:0] arr__U656_out [4:0];
wire arr__U663_clk;
wire [15:0] arr__U663_in [4:0];
wire [15:0] arr__U663_out [4:0];
wire arr__U670_clk;
wire [15:0] arr__U670_in [4:0];
wire [15:0] arr__U670_out [4:0];
wire arr__U677_clk;
wire [15:0] arr__U677_in [4:0];
wire [15:0] arr__U677_out [4:0];
wire arr__U684_clk;
wire [15:0] arr__U684_in [4:0];
wire [15:0] arr__U684_out [4:0];
wire arr__U691_clk;
wire [15:0] arr__U691_in [4:0];
wire [15:0] arr__U691_out [4:0];
wire arr__U698_clk;
wire [15:0] arr__U698_in [4:0];
wire [15:0] arr__U698_out [4:0];
wire arr__U705_clk;
wire [15:0] arr__U705_in [4:0];
wire [15:0] arr__U705_out [4:0];
wire arr__U712_clk;
wire [15:0] arr__U712_in [4:0];
wire [15:0] arr__U712_out [4:0];
wire arr__U719_clk;
wire [15:0] arr__U719_in [4:0];
wire [15:0] arr__U719_out [4:0];
wire arr__U98_clk;
wire [15:0] arr__U98_in [3:0];
wire [15:0] arr__U98_out [3:0];
wire conv_stencil_clk;
wire conv_stencil_flush;
wire conv_stencil_rst_n;
wire conv_stencil_op_hcompute_conv_stencil_1_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_2_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_3_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_4_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire conv_stencil_op_hcompute_conv_stencil_5_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars [4:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire conv_stencil_op_hcompute_conv_stencil_write_wen;
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars [2:0];
wire [15:0] conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire conv_stencil_op_hcompute_hw_output_stencil_read_ren;
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars [3:0];
wire [15:0] conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire delay_reg__U111_clk;
wire delay_reg__U111_in;
wire delay_reg__U111_out;
wire delay_reg__U112_clk;
wire delay_reg__U112_in;
wire delay_reg__U112_out;
wire delay_reg__U159_clk;
wire delay_reg__U159_in;
wire delay_reg__U159_out;
wire delay_reg__U160_clk;
wire delay_reg__U160_in;
wire delay_reg__U160_out;
wire delay_reg__U177_clk;
wire delay_reg__U177_in;
wire delay_reg__U177_out;
wire delay_reg__U178_clk;
wire delay_reg__U178_in;
wire delay_reg__U178_out;
wire delay_reg__U179_clk;
wire delay_reg__U179_in;
wire delay_reg__U179_out;
wire delay_reg__U180_clk;
wire delay_reg__U180_in;
wire delay_reg__U180_out;
wire delay_reg__U181_clk;
wire delay_reg__U181_in;
wire delay_reg__U181_out;
wire delay_reg__U182_clk;
wire delay_reg__U182_in;
wire delay_reg__U182_out;
wire delay_reg__U183_clk;
wire delay_reg__U183_in;
wire delay_reg__U183_out;
wire delay_reg__U184_clk;
wire delay_reg__U184_in;
wire delay_reg__U184_out;
wire delay_reg__U185_clk;
wire delay_reg__U185_in;
wire delay_reg__U185_out;
wire delay_reg__U186_clk;
wire delay_reg__U186_in;
wire delay_reg__U186_out;
wire delay_reg__U187_clk;
wire delay_reg__U187_in;
wire delay_reg__U187_out;
wire delay_reg__U188_clk;
wire delay_reg__U188_in;
wire delay_reg__U188_out;
wire delay_reg__U189_clk;
wire delay_reg__U189_in;
wire delay_reg__U189_out;
wire delay_reg__U190_clk;
wire delay_reg__U190_in;
wire delay_reg__U190_out;
wire delay_reg__U191_clk;
wire delay_reg__U191_in;
wire delay_reg__U191_out;
wire delay_reg__U192_clk;
wire delay_reg__U192_in;
wire delay_reg__U192_out;
wire delay_reg__U193_clk;
wire delay_reg__U193_in;
wire delay_reg__U193_out;
wire delay_reg__U383_clk;
wire delay_reg__U383_in;
wire delay_reg__U383_out;
wire delay_reg__U384_clk;
wire delay_reg__U384_in;
wire delay_reg__U384_out;
wire delay_reg__U401_clk;
wire delay_reg__U401_in;
wire delay_reg__U401_out;
wire delay_reg__U402_clk;
wire delay_reg__U402_in;
wire delay_reg__U402_out;
wire delay_reg__U403_clk;
wire delay_reg__U403_in;
wire delay_reg__U403_out;
wire delay_reg__U404_clk;
wire delay_reg__U404_in;
wire delay_reg__U404_out;
wire delay_reg__U405_clk;
wire delay_reg__U405_in;
wire delay_reg__U405_out;
wire delay_reg__U406_clk;
wire delay_reg__U406_in;
wire delay_reg__U406_out;
wire delay_reg__U407_clk;
wire delay_reg__U407_in;
wire delay_reg__U407_out;
wire delay_reg__U408_clk;
wire delay_reg__U408_in;
wire delay_reg__U408_out;
wire delay_reg__U409_clk;
wire delay_reg__U409_in;
wire delay_reg__U409_out;
wire delay_reg__U410_clk;
wire delay_reg__U410_in;
wire delay_reg__U410_out;
wire delay_reg__U411_clk;
wire delay_reg__U411_in;
wire delay_reg__U411_out;
wire delay_reg__U412_clk;
wire delay_reg__U412_in;
wire delay_reg__U412_out;
wire delay_reg__U413_clk;
wire delay_reg__U413_in;
wire delay_reg__U413_out;
wire delay_reg__U414_clk;
wire delay_reg__U414_in;
wire delay_reg__U414_out;
wire delay_reg__U415_clk;
wire delay_reg__U415_in;
wire delay_reg__U415_out;
wire delay_reg__U416_clk;
wire delay_reg__U416_in;
wire delay_reg__U416_out;
wire delay_reg__U417_clk;
wire delay_reg__U417_in;
wire delay_reg__U417_out;
wire delay_reg__U571_clk;
wire delay_reg__U571_in;
wire delay_reg__U571_out;
wire delay_reg__U572_clk;
wire delay_reg__U572_in;
wire delay_reg__U572_out;
wire delay_reg__U589_clk;
wire delay_reg__U589_in;
wire delay_reg__U589_out;
wire delay_reg__U590_clk;
wire delay_reg__U590_in;
wire delay_reg__U590_out;
wire delay_reg__U591_clk;
wire delay_reg__U591_in;
wire delay_reg__U591_out;
wire delay_reg__U592_clk;
wire delay_reg__U592_in;
wire delay_reg__U592_out;
wire delay_reg__U593_clk;
wire delay_reg__U593_in;
wire delay_reg__U593_out;
wire delay_reg__U594_clk;
wire delay_reg__U594_in;
wire delay_reg__U594_out;
wire delay_reg__U595_clk;
wire delay_reg__U595_in;
wire delay_reg__U595_out;
wire delay_reg__U596_clk;
wire delay_reg__U596_in;
wire delay_reg__U596_out;
wire delay_reg__U597_clk;
wire delay_reg__U597_in;
wire delay_reg__U597_out;
wire delay_reg__U598_clk;
wire delay_reg__U598_in;
wire delay_reg__U598_out;
wire delay_reg__U599_clk;
wire delay_reg__U599_in;
wire delay_reg__U599_out;
wire delay_reg__U600_clk;
wire delay_reg__U600_in;
wire delay_reg__U600_out;
wire delay_reg__U601_clk;
wire delay_reg__U601_in;
wire delay_reg__U601_out;
wire delay_reg__U602_clk;
wire delay_reg__U602_in;
wire delay_reg__U602_out;
wire delay_reg__U603_clk;
wire delay_reg__U603_in;
wire delay_reg__U603_out;
wire delay_reg__U604_clk;
wire delay_reg__U604_in;
wire delay_reg__U604_out;
wire delay_reg__U605_clk;
wire delay_reg__U605_in;
wire delay_reg__U605_out;
wire delay_reg__U95_clk;
wire delay_reg__U95_in;
wire delay_reg__U95_out;
wire delay_reg__U96_clk;
wire delay_reg__U96_in;
wire delay_reg__U96_out;
wire hw_input_global_wrapper_stencil_clk;
wire hw_input_global_wrapper_stencil_flush;
wire hw_input_global_wrapper_stencil_rst_n;
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen;
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars [3:0];
wire [15:0] hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire hw_kernel_global_wrapper_stencil_clk;
wire hw_kernel_global_wrapper_stencil_flush;
wire hw_kernel_global_wrapper_stencil_rst_n;
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen;
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars [4:0];
wire [15:0] hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_conv_stencil_clk;
wire [15:0] op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write [0:0];
wire op_hcompute_conv_stencil_1_clk;
wire [15:0] op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write [0:0];
wire op_hcompute_conv_stencil_1_exe_start_in;
wire op_hcompute_conv_stencil_1_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_port_controller_clk;
wire op_hcompute_conv_stencil_1_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_1_port_controller_d [2:0];
wire op_hcompute_conv_stencil_1_read_start_in;
wire op_hcompute_conv_stencil_1_read_start_out;
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_1_write_start_in;
wire op_hcompute_conv_stencil_1_write_start_out;
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_1_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_clk;
wire [15:0] op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write [0:0];
wire op_hcompute_conv_stencil_2_exe_start_in;
wire op_hcompute_conv_stencil_2_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_port_controller_clk;
wire op_hcompute_conv_stencil_2_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_2_port_controller_d [2:0];
wire op_hcompute_conv_stencil_2_read_start_in;
wire op_hcompute_conv_stencil_2_read_start_out;
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_2_write_start_in;
wire op_hcompute_conv_stencil_2_write_start_out;
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_2_write_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_3_clk;
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read [0:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read [7:0];
wire [15:0] op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write [0:0];
wire op_hcompute_conv_stencil_3_exe_start_in;
wire op_hcompute_conv_stencil_3_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_port_controller_clk;
wire op_hcompute_conv_stencil_3_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_3_port_controller_d [4:0];
wire op_hcompute_conv_stencil_3_read_start_in;
wire op_hcompute_conv_stencil_3_read_start_out;
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_3_write_start_in;
wire op_hcompute_conv_stencil_3_write_start_out;
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_3_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_clk;
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read [0:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read [7:0];
wire [15:0] op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write [0:0];
wire op_hcompute_conv_stencil_4_exe_start_in;
wire op_hcompute_conv_stencil_4_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_port_controller_clk;
wire op_hcompute_conv_stencil_4_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_4_port_controller_d [4:0];
wire op_hcompute_conv_stencil_4_read_start_in;
wire op_hcompute_conv_stencil_4_read_start_out;
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_4_write_start_in;
wire op_hcompute_conv_stencil_4_write_start_out;
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_4_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_clk;
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read [0:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read [7:0];
wire [15:0] op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write [0:0];
wire op_hcompute_conv_stencil_5_exe_start_in;
wire op_hcompute_conv_stencil_5_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_exe_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_port_controller_clk;
wire op_hcompute_conv_stencil_5_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_5_port_controller_d [4:0];
wire op_hcompute_conv_stencil_5_read_start_in;
wire op_hcompute_conv_stencil_5_read_start_out;
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_read_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_5_write_start_in;
wire op_hcompute_conv_stencil_5_write_start_out;
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_conv_stencil_5_write_start_control_vars_out [4:0];
wire op_hcompute_conv_stencil_exe_start_in;
wire op_hcompute_conv_stencil_exe_start_out;
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_exe_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_port_controller_clk;
wire op_hcompute_conv_stencil_port_controller_valid;
wire [15:0] op_hcompute_conv_stencil_port_controller_d [2:0];
wire op_hcompute_conv_stencil_read_start_in;
wire op_hcompute_conv_stencil_read_start_out;
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_read_start_control_vars_out [2:0];
wire op_hcompute_conv_stencil_write_start_in;
wire op_hcompute_conv_stencil_write_start_out;
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_in [2:0];
wire [15:0] op_hcompute_conv_stencil_write_start_control_vars_out [2:0];
wire op_hcompute_hw_input_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_port_controller_d [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out [3:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_clk;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read [0:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write [0:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk;
wire op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out [4:0];
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in;
wire op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in [4:0];
wire [15:0] op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out [4:0];
wire op_hcompute_hw_output_stencil_clk;
wire [15:0] op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read [0:0];
wire [15:0] op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write [0:0];
wire op_hcompute_hw_output_stencil_exe_start_in;
wire op_hcompute_hw_output_stencil_exe_start_out;
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_exe_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_port_controller_clk;
wire op_hcompute_hw_output_stencil_port_controller_valid;
wire [15:0] op_hcompute_hw_output_stencil_port_controller_d [3:0];
wire op_hcompute_hw_output_stencil_read_start_in;
wire op_hcompute_hw_output_stencil_read_start_out;
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_read_start_control_vars_out [3:0];
wire op_hcompute_hw_output_stencil_write_start_in;
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_in [3:0];
wire [15:0] op_hcompute_hw_output_stencil_write_start_control_vars_out [3:0];
assign arr__U104_clk = clk;
assign arr__U104_in[3] = arr__U98_out[3];
assign arr__U104_in[2] = arr__U98_out[2];
assign arr__U104_in[1] = arr__U98_out[1];
assign arr__U104_in[0] = arr__U98_out[0];
array_delay_U105 arr__U104 (
    .clk(arr__U104_clk),
    .in(arr__U104_in),
    .out(arr__U104_out)
);
assign arr__U114_clk = clk;
assign arr__U114_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U114_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U114_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U114_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U115 arr__U114 (
    .clk(arr__U114_clk),
    .in(arr__U114_in),
    .out(arr__U114_out)
);
assign arr__U120_clk = clk;
assign arr__U120_in[3] = arr__U114_out[3];
assign arr__U120_in[2] = arr__U114_out[2];
assign arr__U120_in[1] = arr__U114_out[1];
assign arr__U120_in[0] = arr__U114_out[0];
array_delay_U121 arr__U120 (
    .clk(arr__U120_clk),
    .in(arr__U120_in),
    .out(arr__U120_out)
);
assign arr__U162_clk = clk;
assign arr__U162_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U162_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U162_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U162_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U162_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U163 arr__U162 (
    .clk(arr__U162_clk),
    .in(arr__U162_in),
    .out(arr__U162_out)
);
assign arr__U169_clk = clk;
assign arr__U169_in[4] = arr__U162_out[4];
assign arr__U169_in[3] = arr__U162_out[3];
assign arr__U169_in[2] = arr__U162_out[2];
assign arr__U169_in[1] = arr__U162_out[1];
assign arr__U169_in[0] = arr__U162_out[0];
array_delay_U170 arr__U169 (
    .clk(arr__U169_clk),
    .in(arr__U169_in),
    .out(arr__U169_out)
);
assign arr__U195_clk = clk;
assign arr__U195_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign arr__U195_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign arr__U195_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign arr__U195_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign arr__U195_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
array_delay_U196 arr__U195 (
    .clk(arr__U195_clk),
    .in(arr__U195_in),
    .out(arr__U195_out)
);
assign arr__U202_clk = clk;
assign arr__U202_in[4] = arr__U195_out[4];
assign arr__U202_in[3] = arr__U195_out[3];
assign arr__U202_in[2] = arr__U195_out[2];
assign arr__U202_in[1] = arr__U195_out[1];
assign arr__U202_in[0] = arr__U195_out[0];
array_delay_U203 arr__U202 (
    .clk(arr__U202_clk),
    .in(arr__U202_in),
    .out(arr__U202_out)
);
assign arr__U209_clk = clk;
assign arr__U209_in[4] = arr__U202_out[4];
assign arr__U209_in[3] = arr__U202_out[3];
assign arr__U209_in[2] = arr__U202_out[2];
assign arr__U209_in[1] = arr__U202_out[1];
assign arr__U209_in[0] = arr__U202_out[0];
array_delay_U210 arr__U209 (
    .clk(arr__U209_clk),
    .in(arr__U209_in),
    .out(arr__U209_out)
);
assign arr__U216_clk = clk;
assign arr__U216_in[4] = arr__U209_out[4];
assign arr__U216_in[3] = arr__U209_out[3];
assign arr__U216_in[2] = arr__U209_out[2];
assign arr__U216_in[1] = arr__U209_out[1];
assign arr__U216_in[0] = arr__U209_out[0];
array_delay_U217 arr__U216 (
    .clk(arr__U216_clk),
    .in(arr__U216_in),
    .out(arr__U216_out)
);
assign arr__U223_clk = clk;
assign arr__U223_in[4] = arr__U216_out[4];
assign arr__U223_in[3] = arr__U216_out[3];
assign arr__U223_in[2] = arr__U216_out[2];
assign arr__U223_in[1] = arr__U216_out[1];
assign arr__U223_in[0] = arr__U216_out[0];
array_delay_U224 arr__U223 (
    .clk(arr__U223_clk),
    .in(arr__U223_in),
    .out(arr__U223_out)
);
assign arr__U230_clk = clk;
assign arr__U230_in[4] = arr__U223_out[4];
assign arr__U230_in[3] = arr__U223_out[3];
assign arr__U230_in[2] = arr__U223_out[2];
assign arr__U230_in[1] = arr__U223_out[1];
assign arr__U230_in[0] = arr__U223_out[0];
array_delay_U231 arr__U230 (
    .clk(arr__U230_clk),
    .in(arr__U230_in),
    .out(arr__U230_out)
);
assign arr__U237_clk = clk;
assign arr__U237_in[4] = arr__U230_out[4];
assign arr__U237_in[3] = arr__U230_out[3];
assign arr__U237_in[2] = arr__U230_out[2];
assign arr__U237_in[1] = arr__U230_out[1];
assign arr__U237_in[0] = arr__U230_out[0];
array_delay_U238 arr__U237 (
    .clk(arr__U237_clk),
    .in(arr__U237_in),
    .out(arr__U237_out)
);
assign arr__U244_clk = clk;
assign arr__U244_in[4] = arr__U237_out[4];
assign arr__U244_in[3] = arr__U237_out[3];
assign arr__U244_in[2] = arr__U237_out[2];
assign arr__U244_in[1] = arr__U237_out[1];
assign arr__U244_in[0] = arr__U237_out[0];
array_delay_U245 arr__U244 (
    .clk(arr__U244_clk),
    .in(arr__U244_in),
    .out(arr__U244_out)
);
assign arr__U251_clk = clk;
assign arr__U251_in[4] = arr__U244_out[4];
assign arr__U251_in[3] = arr__U244_out[3];
assign arr__U251_in[2] = arr__U244_out[2];
assign arr__U251_in[1] = arr__U244_out[1];
assign arr__U251_in[0] = arr__U244_out[0];
array_delay_U252 arr__U251 (
    .clk(arr__U251_clk),
    .in(arr__U251_in),
    .out(arr__U251_out)
);
assign arr__U258_clk = clk;
assign arr__U258_in[4] = arr__U251_out[4];
assign arr__U258_in[3] = arr__U251_out[3];
assign arr__U258_in[2] = arr__U251_out[2];
assign arr__U258_in[1] = arr__U251_out[1];
assign arr__U258_in[0] = arr__U251_out[0];
array_delay_U259 arr__U258 (
    .clk(arr__U258_clk),
    .in(arr__U258_in),
    .out(arr__U258_out)
);
assign arr__U265_clk = clk;
assign arr__U265_in[4] = arr__U258_out[4];
assign arr__U265_in[3] = arr__U258_out[3];
assign arr__U265_in[2] = arr__U258_out[2];
assign arr__U265_in[1] = arr__U258_out[1];
assign arr__U265_in[0] = arr__U258_out[0];
array_delay_U266 arr__U265 (
    .clk(arr__U265_clk),
    .in(arr__U265_in),
    .out(arr__U265_out)
);
assign arr__U272_clk = clk;
assign arr__U272_in[4] = arr__U265_out[4];
assign arr__U272_in[3] = arr__U265_out[3];
assign arr__U272_in[2] = arr__U265_out[2];
assign arr__U272_in[1] = arr__U265_out[1];
assign arr__U272_in[0] = arr__U265_out[0];
array_delay_U273 arr__U272 (
    .clk(arr__U272_clk),
    .in(arr__U272_in),
    .out(arr__U272_out)
);
assign arr__U279_clk = clk;
assign arr__U279_in[4] = arr__U272_out[4];
assign arr__U279_in[3] = arr__U272_out[3];
assign arr__U279_in[2] = arr__U272_out[2];
assign arr__U279_in[1] = arr__U272_out[1];
assign arr__U279_in[0] = arr__U272_out[0];
array_delay_U280 arr__U279 (
    .clk(arr__U279_clk),
    .in(arr__U279_in),
    .out(arr__U279_out)
);
assign arr__U286_clk = clk;
assign arr__U286_in[4] = arr__U279_out[4];
assign arr__U286_in[3] = arr__U279_out[3];
assign arr__U286_in[2] = arr__U279_out[2];
assign arr__U286_in[1] = arr__U279_out[1];
assign arr__U286_in[0] = arr__U279_out[0];
array_delay_U287 arr__U286 (
    .clk(arr__U286_clk),
    .in(arr__U286_in),
    .out(arr__U286_out)
);
assign arr__U293_clk = clk;
assign arr__U293_in[4] = arr__U286_out[4];
assign arr__U293_in[3] = arr__U286_out[3];
assign arr__U293_in[2] = arr__U286_out[2];
assign arr__U293_in[1] = arr__U286_out[1];
assign arr__U293_in[0] = arr__U286_out[0];
array_delay_U294 arr__U293 (
    .clk(arr__U293_clk),
    .in(arr__U293_in),
    .out(arr__U293_out)
);
assign arr__U300_clk = clk;
assign arr__U300_in[4] = arr__U293_out[4];
assign arr__U300_in[3] = arr__U293_out[3];
assign arr__U300_in[2] = arr__U293_out[2];
assign arr__U300_in[1] = arr__U293_out[1];
assign arr__U300_in[0] = arr__U293_out[0];
array_delay_U301 arr__U300 (
    .clk(arr__U300_clk),
    .in(arr__U300_in),
    .out(arr__U300_out)
);
assign arr__U307_clk = clk;
assign arr__U307_in[4] = arr__U300_out[4];
assign arr__U307_in[3] = arr__U300_out[3];
assign arr__U307_in[2] = arr__U300_out[2];
assign arr__U307_in[1] = arr__U300_out[1];
assign arr__U307_in[0] = arr__U300_out[0];
array_delay_U308 arr__U307 (
    .clk(arr__U307_clk),
    .in(arr__U307_in),
    .out(arr__U307_out)
);
assign arr__U386_clk = clk;
assign arr__U386_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U386_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U386_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U386_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U386_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U387 arr__U386 (
    .clk(arr__U386_clk),
    .in(arr__U386_in),
    .out(arr__U386_out)
);
assign arr__U393_clk = clk;
assign arr__U393_in[4] = arr__U386_out[4];
assign arr__U393_in[3] = arr__U386_out[3];
assign arr__U393_in[2] = arr__U386_out[2];
assign arr__U393_in[1] = arr__U386_out[1];
assign arr__U393_in[0] = arr__U386_out[0];
array_delay_U394 arr__U393 (
    .clk(arr__U393_clk),
    .in(arr__U393_in),
    .out(arr__U393_out)
);
assign arr__U419_clk = clk;
assign arr__U419_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign arr__U419_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign arr__U419_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign arr__U419_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign arr__U419_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
array_delay_U420 arr__U419 (
    .clk(arr__U419_clk),
    .in(arr__U419_in),
    .out(arr__U419_out)
);
assign arr__U426_clk = clk;
assign arr__U426_in[4] = arr__U419_out[4];
assign arr__U426_in[3] = arr__U419_out[3];
assign arr__U426_in[2] = arr__U419_out[2];
assign arr__U426_in[1] = arr__U419_out[1];
assign arr__U426_in[0] = arr__U419_out[0];
array_delay_U427 arr__U426 (
    .clk(arr__U426_clk),
    .in(arr__U426_in),
    .out(arr__U426_out)
);
assign arr__U433_clk = clk;
assign arr__U433_in[4] = arr__U426_out[4];
assign arr__U433_in[3] = arr__U426_out[3];
assign arr__U433_in[2] = arr__U426_out[2];
assign arr__U433_in[1] = arr__U426_out[1];
assign arr__U433_in[0] = arr__U426_out[0];
array_delay_U434 arr__U433 (
    .clk(arr__U433_clk),
    .in(arr__U433_in),
    .out(arr__U433_out)
);
assign arr__U440_clk = clk;
assign arr__U440_in[4] = arr__U433_out[4];
assign arr__U440_in[3] = arr__U433_out[3];
assign arr__U440_in[2] = arr__U433_out[2];
assign arr__U440_in[1] = arr__U433_out[1];
assign arr__U440_in[0] = arr__U433_out[0];
array_delay_U441 arr__U440 (
    .clk(arr__U440_clk),
    .in(arr__U440_in),
    .out(arr__U440_out)
);
assign arr__U447_clk = clk;
assign arr__U447_in[4] = arr__U440_out[4];
assign arr__U447_in[3] = arr__U440_out[3];
assign arr__U447_in[2] = arr__U440_out[2];
assign arr__U447_in[1] = arr__U440_out[1];
assign arr__U447_in[0] = arr__U440_out[0];
array_delay_U448 arr__U447 (
    .clk(arr__U447_clk),
    .in(arr__U447_in),
    .out(arr__U447_out)
);
assign arr__U454_clk = clk;
assign arr__U454_in[4] = arr__U447_out[4];
assign arr__U454_in[3] = arr__U447_out[3];
assign arr__U454_in[2] = arr__U447_out[2];
assign arr__U454_in[1] = arr__U447_out[1];
assign arr__U454_in[0] = arr__U447_out[0];
array_delay_U455 arr__U454 (
    .clk(arr__U454_clk),
    .in(arr__U454_in),
    .out(arr__U454_out)
);
assign arr__U461_clk = clk;
assign arr__U461_in[4] = arr__U454_out[4];
assign arr__U461_in[3] = arr__U454_out[3];
assign arr__U461_in[2] = arr__U454_out[2];
assign arr__U461_in[1] = arr__U454_out[1];
assign arr__U461_in[0] = arr__U454_out[0];
array_delay_U462 arr__U461 (
    .clk(arr__U461_clk),
    .in(arr__U461_in),
    .out(arr__U461_out)
);
assign arr__U468_clk = clk;
assign arr__U468_in[4] = arr__U461_out[4];
assign arr__U468_in[3] = arr__U461_out[3];
assign arr__U468_in[2] = arr__U461_out[2];
assign arr__U468_in[1] = arr__U461_out[1];
assign arr__U468_in[0] = arr__U461_out[0];
array_delay_U469 arr__U468 (
    .clk(arr__U468_clk),
    .in(arr__U468_in),
    .out(arr__U468_out)
);
assign arr__U475_clk = clk;
assign arr__U475_in[4] = arr__U468_out[4];
assign arr__U475_in[3] = arr__U468_out[3];
assign arr__U475_in[2] = arr__U468_out[2];
assign arr__U475_in[1] = arr__U468_out[1];
assign arr__U475_in[0] = arr__U468_out[0];
array_delay_U476 arr__U475 (
    .clk(arr__U475_clk),
    .in(arr__U475_in),
    .out(arr__U475_out)
);
assign arr__U482_clk = clk;
assign arr__U482_in[4] = arr__U475_out[4];
assign arr__U482_in[3] = arr__U475_out[3];
assign arr__U482_in[2] = arr__U475_out[2];
assign arr__U482_in[1] = arr__U475_out[1];
assign arr__U482_in[0] = arr__U475_out[0];
array_delay_U483 arr__U482 (
    .clk(arr__U482_clk),
    .in(arr__U482_in),
    .out(arr__U482_out)
);
assign arr__U489_clk = clk;
assign arr__U489_in[4] = arr__U482_out[4];
assign arr__U489_in[3] = arr__U482_out[3];
assign arr__U489_in[2] = arr__U482_out[2];
assign arr__U489_in[1] = arr__U482_out[1];
assign arr__U489_in[0] = arr__U482_out[0];
array_delay_U490 arr__U489 (
    .clk(arr__U489_clk),
    .in(arr__U489_in),
    .out(arr__U489_out)
);
assign arr__U496_clk = clk;
assign arr__U496_in[4] = arr__U489_out[4];
assign arr__U496_in[3] = arr__U489_out[3];
assign arr__U496_in[2] = arr__U489_out[2];
assign arr__U496_in[1] = arr__U489_out[1];
assign arr__U496_in[0] = arr__U489_out[0];
array_delay_U497 arr__U496 (
    .clk(arr__U496_clk),
    .in(arr__U496_in),
    .out(arr__U496_out)
);
assign arr__U503_clk = clk;
assign arr__U503_in[4] = arr__U496_out[4];
assign arr__U503_in[3] = arr__U496_out[3];
assign arr__U503_in[2] = arr__U496_out[2];
assign arr__U503_in[1] = arr__U496_out[1];
assign arr__U503_in[0] = arr__U496_out[0];
array_delay_U504 arr__U503 (
    .clk(arr__U503_clk),
    .in(arr__U503_in),
    .out(arr__U503_out)
);
assign arr__U510_clk = clk;
assign arr__U510_in[4] = arr__U503_out[4];
assign arr__U510_in[3] = arr__U503_out[3];
assign arr__U510_in[2] = arr__U503_out[2];
assign arr__U510_in[1] = arr__U503_out[1];
assign arr__U510_in[0] = arr__U503_out[0];
array_delay_U511 arr__U510 (
    .clk(arr__U510_clk),
    .in(arr__U510_in),
    .out(arr__U510_out)
);
assign arr__U517_clk = clk;
assign arr__U517_in[4] = arr__U510_out[4];
assign arr__U517_in[3] = arr__U510_out[3];
assign arr__U517_in[2] = arr__U510_out[2];
assign arr__U517_in[1] = arr__U510_out[1];
assign arr__U517_in[0] = arr__U510_out[0];
array_delay_U518 arr__U517 (
    .clk(arr__U517_clk),
    .in(arr__U517_in),
    .out(arr__U517_out)
);
assign arr__U524_clk = clk;
assign arr__U524_in[4] = arr__U517_out[4];
assign arr__U524_in[3] = arr__U517_out[3];
assign arr__U524_in[2] = arr__U517_out[2];
assign arr__U524_in[1] = arr__U517_out[1];
assign arr__U524_in[0] = arr__U517_out[0];
array_delay_U525 arr__U524 (
    .clk(arr__U524_clk),
    .in(arr__U524_in),
    .out(arr__U524_out)
);
assign arr__U531_clk = clk;
assign arr__U531_in[4] = arr__U524_out[4];
assign arr__U531_in[3] = arr__U524_out[3];
assign arr__U531_in[2] = arr__U524_out[2];
assign arr__U531_in[1] = arr__U524_out[1];
assign arr__U531_in[0] = arr__U524_out[0];
array_delay_U532 arr__U531 (
    .clk(arr__U531_clk),
    .in(arr__U531_in),
    .out(arr__U531_out)
);
assign arr__U574_clk = clk;
assign arr__U574_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U574_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U574_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U574_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U574_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U575 arr__U574 (
    .clk(arr__U574_clk),
    .in(arr__U574_in),
    .out(arr__U574_out)
);
assign arr__U581_clk = clk;
assign arr__U581_in[4] = arr__U574_out[4];
assign arr__U581_in[3] = arr__U574_out[3];
assign arr__U581_in[2] = arr__U574_out[2];
assign arr__U581_in[1] = arr__U574_out[1];
assign arr__U581_in[0] = arr__U574_out[0];
array_delay_U582 arr__U581 (
    .clk(arr__U581_clk),
    .in(arr__U581_in),
    .out(arr__U581_out)
);
assign arr__U607_clk = clk;
assign arr__U607_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign arr__U607_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign arr__U607_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign arr__U607_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign arr__U607_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
array_delay_U608 arr__U607 (
    .clk(arr__U607_clk),
    .in(arr__U607_in),
    .out(arr__U607_out)
);
assign arr__U614_clk = clk;
assign arr__U614_in[4] = arr__U607_out[4];
assign arr__U614_in[3] = arr__U607_out[3];
assign arr__U614_in[2] = arr__U607_out[2];
assign arr__U614_in[1] = arr__U607_out[1];
assign arr__U614_in[0] = arr__U607_out[0];
array_delay_U615 arr__U614 (
    .clk(arr__U614_clk),
    .in(arr__U614_in),
    .out(arr__U614_out)
);
assign arr__U621_clk = clk;
assign arr__U621_in[4] = arr__U614_out[4];
assign arr__U621_in[3] = arr__U614_out[3];
assign arr__U621_in[2] = arr__U614_out[2];
assign arr__U621_in[1] = arr__U614_out[1];
assign arr__U621_in[0] = arr__U614_out[0];
array_delay_U622 arr__U621 (
    .clk(arr__U621_clk),
    .in(arr__U621_in),
    .out(arr__U621_out)
);
assign arr__U628_clk = clk;
assign arr__U628_in[4] = arr__U621_out[4];
assign arr__U628_in[3] = arr__U621_out[3];
assign arr__U628_in[2] = arr__U621_out[2];
assign arr__U628_in[1] = arr__U621_out[1];
assign arr__U628_in[0] = arr__U621_out[0];
array_delay_U629 arr__U628 (
    .clk(arr__U628_clk),
    .in(arr__U628_in),
    .out(arr__U628_out)
);
assign arr__U635_clk = clk;
assign arr__U635_in[4] = arr__U628_out[4];
assign arr__U635_in[3] = arr__U628_out[3];
assign arr__U635_in[2] = arr__U628_out[2];
assign arr__U635_in[1] = arr__U628_out[1];
assign arr__U635_in[0] = arr__U628_out[0];
array_delay_U636 arr__U635 (
    .clk(arr__U635_clk),
    .in(arr__U635_in),
    .out(arr__U635_out)
);
assign arr__U642_clk = clk;
assign arr__U642_in[4] = arr__U635_out[4];
assign arr__U642_in[3] = arr__U635_out[3];
assign arr__U642_in[2] = arr__U635_out[2];
assign arr__U642_in[1] = arr__U635_out[1];
assign arr__U642_in[0] = arr__U635_out[0];
array_delay_U643 arr__U642 (
    .clk(arr__U642_clk),
    .in(arr__U642_in),
    .out(arr__U642_out)
);
assign arr__U649_clk = clk;
assign arr__U649_in[4] = arr__U642_out[4];
assign arr__U649_in[3] = arr__U642_out[3];
assign arr__U649_in[2] = arr__U642_out[2];
assign arr__U649_in[1] = arr__U642_out[1];
assign arr__U649_in[0] = arr__U642_out[0];
array_delay_U650 arr__U649 (
    .clk(arr__U649_clk),
    .in(arr__U649_in),
    .out(arr__U649_out)
);
assign arr__U656_clk = clk;
assign arr__U656_in[4] = arr__U649_out[4];
assign arr__U656_in[3] = arr__U649_out[3];
assign arr__U656_in[2] = arr__U649_out[2];
assign arr__U656_in[1] = arr__U649_out[1];
assign arr__U656_in[0] = arr__U649_out[0];
array_delay_U657 arr__U656 (
    .clk(arr__U656_clk),
    .in(arr__U656_in),
    .out(arr__U656_out)
);
assign arr__U663_clk = clk;
assign arr__U663_in[4] = arr__U656_out[4];
assign arr__U663_in[3] = arr__U656_out[3];
assign arr__U663_in[2] = arr__U656_out[2];
assign arr__U663_in[1] = arr__U656_out[1];
assign arr__U663_in[0] = arr__U656_out[0];
array_delay_U664 arr__U663 (
    .clk(arr__U663_clk),
    .in(arr__U663_in),
    .out(arr__U663_out)
);
assign arr__U670_clk = clk;
assign arr__U670_in[4] = arr__U663_out[4];
assign arr__U670_in[3] = arr__U663_out[3];
assign arr__U670_in[2] = arr__U663_out[2];
assign arr__U670_in[1] = arr__U663_out[1];
assign arr__U670_in[0] = arr__U663_out[0];
array_delay_U671 arr__U670 (
    .clk(arr__U670_clk),
    .in(arr__U670_in),
    .out(arr__U670_out)
);
assign arr__U677_clk = clk;
assign arr__U677_in[4] = arr__U670_out[4];
assign arr__U677_in[3] = arr__U670_out[3];
assign arr__U677_in[2] = arr__U670_out[2];
assign arr__U677_in[1] = arr__U670_out[1];
assign arr__U677_in[0] = arr__U670_out[0];
array_delay_U678 arr__U677 (
    .clk(arr__U677_clk),
    .in(arr__U677_in),
    .out(arr__U677_out)
);
assign arr__U684_clk = clk;
assign arr__U684_in[4] = arr__U677_out[4];
assign arr__U684_in[3] = arr__U677_out[3];
assign arr__U684_in[2] = arr__U677_out[2];
assign arr__U684_in[1] = arr__U677_out[1];
assign arr__U684_in[0] = arr__U677_out[0];
array_delay_U685 arr__U684 (
    .clk(arr__U684_clk),
    .in(arr__U684_in),
    .out(arr__U684_out)
);
assign arr__U691_clk = clk;
assign arr__U691_in[4] = arr__U684_out[4];
assign arr__U691_in[3] = arr__U684_out[3];
assign arr__U691_in[2] = arr__U684_out[2];
assign arr__U691_in[1] = arr__U684_out[1];
assign arr__U691_in[0] = arr__U684_out[0];
array_delay_U692 arr__U691 (
    .clk(arr__U691_clk),
    .in(arr__U691_in),
    .out(arr__U691_out)
);
assign arr__U698_clk = clk;
assign arr__U698_in[4] = arr__U691_out[4];
assign arr__U698_in[3] = arr__U691_out[3];
assign arr__U698_in[2] = arr__U691_out[2];
assign arr__U698_in[1] = arr__U691_out[1];
assign arr__U698_in[0] = arr__U691_out[0];
array_delay_U699 arr__U698 (
    .clk(arr__U698_clk),
    .in(arr__U698_in),
    .out(arr__U698_out)
);
assign arr__U705_clk = clk;
assign arr__U705_in[4] = arr__U698_out[4];
assign arr__U705_in[3] = arr__U698_out[3];
assign arr__U705_in[2] = arr__U698_out[2];
assign arr__U705_in[1] = arr__U698_out[1];
assign arr__U705_in[0] = arr__U698_out[0];
array_delay_U706 arr__U705 (
    .clk(arr__U705_clk),
    .in(arr__U705_in),
    .out(arr__U705_out)
);
assign arr__U712_clk = clk;
assign arr__U712_in[4] = arr__U705_out[4];
assign arr__U712_in[3] = arr__U705_out[3];
assign arr__U712_in[2] = arr__U705_out[2];
assign arr__U712_in[1] = arr__U705_out[1];
assign arr__U712_in[0] = arr__U705_out[0];
array_delay_U713 arr__U712 (
    .clk(arr__U712_clk),
    .in(arr__U712_in),
    .out(arr__U712_out)
);
assign arr__U719_clk = clk;
assign arr__U719_in[4] = arr__U712_out[4];
assign arr__U719_in[3] = arr__U712_out[3];
assign arr__U719_in[2] = arr__U712_out[2];
assign arr__U719_in[1] = arr__U712_out[1];
assign arr__U719_in[0] = arr__U712_out[0];
array_delay_U720 arr__U719 (
    .clk(arr__U719_clk),
    .in(arr__U719_in),
    .out(arr__U719_out)
);
assign arr__U98_clk = clk;
assign arr__U98_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign arr__U98_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign arr__U98_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign arr__U98_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
array_delay_U99 arr__U98 (
    .clk(arr__U98_clk),
    .in(arr__U98_in),
    .out(arr__U98_out)
);
assign conv_stencil_clk = clk;
assign conv_stencil_flush = flush;
assign conv_stencil_rst_n = rst_n;
assign conv_stencil_op_hcompute_conv_stencil_1_write_wen = op_hcompute_conv_stencil_1_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[2] = op_hcompute_conv_stencil_1_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[1] = op_hcompute_conv_stencil_1_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars[0] = op_hcompute_conv_stencil_1_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_1_write[0] = op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write_wen = op_hcompute_conv_stencil_2_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[2] = op_hcompute_conv_stencil_2_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[1] = op_hcompute_conv_stencil_2_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars[0] = op_hcompute_conv_stencil_2_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_2_write[0] = op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write[0];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write_wen = op_hcompute_conv_stencil_3_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[4] = op_hcompute_conv_stencil_3_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[3] = op_hcompute_conv_stencil_3_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[2] = op_hcompute_conv_stencil_3_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[1] = op_hcompute_conv_stencil_3_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars[0] = op_hcompute_conv_stencil_3_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_3_write[0] = op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write[0];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write_wen = op_hcompute_conv_stencil_4_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[4] = op_hcompute_conv_stencil_4_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[3] = op_hcompute_conv_stencil_4_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[2] = op_hcompute_conv_stencil_4_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[1] = op_hcompute_conv_stencil_4_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars[0] = op_hcompute_conv_stencil_4_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_4_write[0] = op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write[0];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write_wen = op_hcompute_conv_stencil_5_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[4] = op_hcompute_conv_stencil_5_write_start_control_vars_out[4];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[3] = op_hcompute_conv_stencil_5_write_start_control_vars_out[3];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[2] = op_hcompute_conv_stencil_5_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[1] = op_hcompute_conv_stencil_5_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars[0] = op_hcompute_conv_stencil_5_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_5_write[0] = op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write[0];
assign conv_stencil_op_hcompute_conv_stencil_write_wen = op_hcompute_conv_stencil_write_start_out;
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[2] = op_hcompute_conv_stencil_write_start_control_vars_out[2];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[1] = op_hcompute_conv_stencil_write_start_control_vars_out[1];
assign conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars[0] = op_hcompute_conv_stencil_write_start_control_vars_out[0];
assign conv_stencil_op_hcompute_conv_stencil_write[0] = op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write[0];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ren = op_hcompute_hw_output_stencil_read_start_out;
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
conv_stencil_ub conv_stencil (
    .clk(conv_stencil_clk),
    .flush(conv_stencil_flush),
    .rst_n(conv_stencil_rst_n),
    .op_hcompute_conv_stencil_1_write_wen(conv_stencil_op_hcompute_conv_stencil_1_write_wen),
    .op_hcompute_conv_stencil_1_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_1_write_ctrl_vars),
    .op_hcompute_conv_stencil_1_write(conv_stencil_op_hcompute_conv_stencil_1_write),
    .op_hcompute_conv_stencil_2_write_wen(conv_stencil_op_hcompute_conv_stencil_2_write_wen),
    .op_hcompute_conv_stencil_2_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_2_write_ctrl_vars),
    .op_hcompute_conv_stencil_2_write(conv_stencil_op_hcompute_conv_stencil_2_write),
    .op_hcompute_conv_stencil_3_read_ren(conv_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(conv_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_3_write_wen(conv_stencil_op_hcompute_conv_stencil_3_write_wen),
    .op_hcompute_conv_stencil_3_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_3_write_ctrl_vars),
    .op_hcompute_conv_stencil_3_write(conv_stencil_op_hcompute_conv_stencil_3_write),
    .op_hcompute_conv_stencil_4_read_ren(conv_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(conv_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_4_write_wen(conv_stencil_op_hcompute_conv_stencil_4_write_wen),
    .op_hcompute_conv_stencil_4_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_4_write_ctrl_vars),
    .op_hcompute_conv_stencil_4_write(conv_stencil_op_hcompute_conv_stencil_4_write),
    .op_hcompute_conv_stencil_5_read_ren(conv_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(conv_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_conv_stencil_5_write_wen(conv_stencil_op_hcompute_conv_stencil_5_write_wen),
    .op_hcompute_conv_stencil_5_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_5_write_ctrl_vars),
    .op_hcompute_conv_stencil_5_write(conv_stencil_op_hcompute_conv_stencil_5_write),
    .op_hcompute_conv_stencil_write_wen(conv_stencil_op_hcompute_conv_stencil_write_wen),
    .op_hcompute_conv_stencil_write_ctrl_vars(conv_stencil_op_hcompute_conv_stencil_write_ctrl_vars),
    .op_hcompute_conv_stencil_write(conv_stencil_op_hcompute_conv_stencil_write),
    .op_hcompute_hw_output_stencil_read_ren(conv_stencil_op_hcompute_hw_output_stencil_read_ren),
    .op_hcompute_hw_output_stencil_read_ctrl_vars(conv_stencil_op_hcompute_hw_output_stencil_read_ctrl_vars),
    .op_hcompute_hw_output_stencil_read(conv_stencil_op_hcompute_hw_output_stencil_read)
);
assign delay_reg__U111_clk = clk;
assign delay_reg__U111_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U111 (
    .clk(delay_reg__U111_clk),
    .in(delay_reg__U111_in),
    .out(delay_reg__U111_out)
);
assign delay_reg__U112_clk = clk;
assign delay_reg__U112_in = delay_reg__U111_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U112 (
    .clk(delay_reg__U112_clk),
    .in(delay_reg__U112_in),
    .out(delay_reg__U112_out)
);
assign delay_reg__U159_clk = clk;
assign delay_reg__U159_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U159 (
    .clk(delay_reg__U159_clk),
    .in(delay_reg__U159_in),
    .out(delay_reg__U159_out)
);
assign delay_reg__U160_clk = clk;
assign delay_reg__U160_in = delay_reg__U159_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U160 (
    .clk(delay_reg__U160_clk),
    .in(delay_reg__U160_in),
    .out(delay_reg__U160_out)
);
assign delay_reg__U177_clk = clk;
assign delay_reg__U177_in = op_hcompute_conv_stencil_5_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U177 (
    .clk(delay_reg__U177_clk),
    .in(delay_reg__U177_in),
    .out(delay_reg__U177_out)
);
assign delay_reg__U178_clk = clk;
assign delay_reg__U178_in = delay_reg__U177_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U178 (
    .clk(delay_reg__U178_clk),
    .in(delay_reg__U178_in),
    .out(delay_reg__U178_out)
);
assign delay_reg__U179_clk = clk;
assign delay_reg__U179_in = delay_reg__U178_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U179 (
    .clk(delay_reg__U179_clk),
    .in(delay_reg__U179_in),
    .out(delay_reg__U179_out)
);
assign delay_reg__U180_clk = clk;
assign delay_reg__U180_in = delay_reg__U179_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U180 (
    .clk(delay_reg__U180_clk),
    .in(delay_reg__U180_in),
    .out(delay_reg__U180_out)
);
assign delay_reg__U181_clk = clk;
assign delay_reg__U181_in = delay_reg__U180_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U181 (
    .clk(delay_reg__U181_clk),
    .in(delay_reg__U181_in),
    .out(delay_reg__U181_out)
);
assign delay_reg__U182_clk = clk;
assign delay_reg__U182_in = delay_reg__U181_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U182 (
    .clk(delay_reg__U182_clk),
    .in(delay_reg__U182_in),
    .out(delay_reg__U182_out)
);
assign delay_reg__U183_clk = clk;
assign delay_reg__U183_in = delay_reg__U182_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U183 (
    .clk(delay_reg__U183_clk),
    .in(delay_reg__U183_in),
    .out(delay_reg__U183_out)
);
assign delay_reg__U184_clk = clk;
assign delay_reg__U184_in = delay_reg__U183_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U184 (
    .clk(delay_reg__U184_clk),
    .in(delay_reg__U184_in),
    .out(delay_reg__U184_out)
);
assign delay_reg__U185_clk = clk;
assign delay_reg__U185_in = delay_reg__U184_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U185 (
    .clk(delay_reg__U185_clk),
    .in(delay_reg__U185_in),
    .out(delay_reg__U185_out)
);
assign delay_reg__U186_clk = clk;
assign delay_reg__U186_in = delay_reg__U185_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U186 (
    .clk(delay_reg__U186_clk),
    .in(delay_reg__U186_in),
    .out(delay_reg__U186_out)
);
assign delay_reg__U187_clk = clk;
assign delay_reg__U187_in = delay_reg__U186_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U187 (
    .clk(delay_reg__U187_clk),
    .in(delay_reg__U187_in),
    .out(delay_reg__U187_out)
);
assign delay_reg__U188_clk = clk;
assign delay_reg__U188_in = delay_reg__U187_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U188 (
    .clk(delay_reg__U188_clk),
    .in(delay_reg__U188_in),
    .out(delay_reg__U188_out)
);
assign delay_reg__U189_clk = clk;
assign delay_reg__U189_in = delay_reg__U188_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U189 (
    .clk(delay_reg__U189_clk),
    .in(delay_reg__U189_in),
    .out(delay_reg__U189_out)
);
assign delay_reg__U190_clk = clk;
assign delay_reg__U190_in = delay_reg__U189_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U190 (
    .clk(delay_reg__U190_clk),
    .in(delay_reg__U190_in),
    .out(delay_reg__U190_out)
);
assign delay_reg__U191_clk = clk;
assign delay_reg__U191_in = delay_reg__U190_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U191 (
    .clk(delay_reg__U191_clk),
    .in(delay_reg__U191_in),
    .out(delay_reg__U191_out)
);
assign delay_reg__U192_clk = clk;
assign delay_reg__U192_in = delay_reg__U191_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U192 (
    .clk(delay_reg__U192_clk),
    .in(delay_reg__U192_in),
    .out(delay_reg__U192_out)
);
assign delay_reg__U193_clk = clk;
assign delay_reg__U193_in = delay_reg__U192_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U193 (
    .clk(delay_reg__U193_clk),
    .in(delay_reg__U193_in),
    .out(delay_reg__U193_out)
);
assign delay_reg__U383_clk = clk;
assign delay_reg__U383_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U383 (
    .clk(delay_reg__U383_clk),
    .in(delay_reg__U383_in),
    .out(delay_reg__U383_out)
);
assign delay_reg__U384_clk = clk;
assign delay_reg__U384_in = delay_reg__U383_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U384 (
    .clk(delay_reg__U384_clk),
    .in(delay_reg__U384_in),
    .out(delay_reg__U384_out)
);
assign delay_reg__U401_clk = clk;
assign delay_reg__U401_in = op_hcompute_conv_stencil_4_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U401 (
    .clk(delay_reg__U401_clk),
    .in(delay_reg__U401_in),
    .out(delay_reg__U401_out)
);
assign delay_reg__U402_clk = clk;
assign delay_reg__U402_in = delay_reg__U401_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U402 (
    .clk(delay_reg__U402_clk),
    .in(delay_reg__U402_in),
    .out(delay_reg__U402_out)
);
assign delay_reg__U403_clk = clk;
assign delay_reg__U403_in = delay_reg__U402_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U403 (
    .clk(delay_reg__U403_clk),
    .in(delay_reg__U403_in),
    .out(delay_reg__U403_out)
);
assign delay_reg__U404_clk = clk;
assign delay_reg__U404_in = delay_reg__U403_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U404 (
    .clk(delay_reg__U404_clk),
    .in(delay_reg__U404_in),
    .out(delay_reg__U404_out)
);
assign delay_reg__U405_clk = clk;
assign delay_reg__U405_in = delay_reg__U404_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U405 (
    .clk(delay_reg__U405_clk),
    .in(delay_reg__U405_in),
    .out(delay_reg__U405_out)
);
assign delay_reg__U406_clk = clk;
assign delay_reg__U406_in = delay_reg__U405_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U406 (
    .clk(delay_reg__U406_clk),
    .in(delay_reg__U406_in),
    .out(delay_reg__U406_out)
);
assign delay_reg__U407_clk = clk;
assign delay_reg__U407_in = delay_reg__U406_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U407 (
    .clk(delay_reg__U407_clk),
    .in(delay_reg__U407_in),
    .out(delay_reg__U407_out)
);
assign delay_reg__U408_clk = clk;
assign delay_reg__U408_in = delay_reg__U407_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U408 (
    .clk(delay_reg__U408_clk),
    .in(delay_reg__U408_in),
    .out(delay_reg__U408_out)
);
assign delay_reg__U409_clk = clk;
assign delay_reg__U409_in = delay_reg__U408_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U409 (
    .clk(delay_reg__U409_clk),
    .in(delay_reg__U409_in),
    .out(delay_reg__U409_out)
);
assign delay_reg__U410_clk = clk;
assign delay_reg__U410_in = delay_reg__U409_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U410 (
    .clk(delay_reg__U410_clk),
    .in(delay_reg__U410_in),
    .out(delay_reg__U410_out)
);
assign delay_reg__U411_clk = clk;
assign delay_reg__U411_in = delay_reg__U410_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U411 (
    .clk(delay_reg__U411_clk),
    .in(delay_reg__U411_in),
    .out(delay_reg__U411_out)
);
assign delay_reg__U412_clk = clk;
assign delay_reg__U412_in = delay_reg__U411_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U412 (
    .clk(delay_reg__U412_clk),
    .in(delay_reg__U412_in),
    .out(delay_reg__U412_out)
);
assign delay_reg__U413_clk = clk;
assign delay_reg__U413_in = delay_reg__U412_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U413 (
    .clk(delay_reg__U413_clk),
    .in(delay_reg__U413_in),
    .out(delay_reg__U413_out)
);
assign delay_reg__U414_clk = clk;
assign delay_reg__U414_in = delay_reg__U413_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U414 (
    .clk(delay_reg__U414_clk),
    .in(delay_reg__U414_in),
    .out(delay_reg__U414_out)
);
assign delay_reg__U415_clk = clk;
assign delay_reg__U415_in = delay_reg__U414_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U415 (
    .clk(delay_reg__U415_clk),
    .in(delay_reg__U415_in),
    .out(delay_reg__U415_out)
);
assign delay_reg__U416_clk = clk;
assign delay_reg__U416_in = delay_reg__U415_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U416 (
    .clk(delay_reg__U416_clk),
    .in(delay_reg__U416_in),
    .out(delay_reg__U416_out)
);
assign delay_reg__U417_clk = clk;
assign delay_reg__U417_in = delay_reg__U416_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U417 (
    .clk(delay_reg__U417_clk),
    .in(delay_reg__U417_in),
    .out(delay_reg__U417_out)
);
assign delay_reg__U571_clk = clk;
assign delay_reg__U571_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U571 (
    .clk(delay_reg__U571_clk),
    .in(delay_reg__U571_in),
    .out(delay_reg__U571_out)
);
assign delay_reg__U572_clk = clk;
assign delay_reg__U572_in = delay_reg__U571_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U572 (
    .clk(delay_reg__U572_clk),
    .in(delay_reg__U572_in),
    .out(delay_reg__U572_out)
);
assign delay_reg__U589_clk = clk;
assign delay_reg__U589_in = op_hcompute_conv_stencil_3_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U589 (
    .clk(delay_reg__U589_clk),
    .in(delay_reg__U589_in),
    .out(delay_reg__U589_out)
);
assign delay_reg__U590_clk = clk;
assign delay_reg__U590_in = delay_reg__U589_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U590 (
    .clk(delay_reg__U590_clk),
    .in(delay_reg__U590_in),
    .out(delay_reg__U590_out)
);
assign delay_reg__U591_clk = clk;
assign delay_reg__U591_in = delay_reg__U590_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U591 (
    .clk(delay_reg__U591_clk),
    .in(delay_reg__U591_in),
    .out(delay_reg__U591_out)
);
assign delay_reg__U592_clk = clk;
assign delay_reg__U592_in = delay_reg__U591_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U592 (
    .clk(delay_reg__U592_clk),
    .in(delay_reg__U592_in),
    .out(delay_reg__U592_out)
);
assign delay_reg__U593_clk = clk;
assign delay_reg__U593_in = delay_reg__U592_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U593 (
    .clk(delay_reg__U593_clk),
    .in(delay_reg__U593_in),
    .out(delay_reg__U593_out)
);
assign delay_reg__U594_clk = clk;
assign delay_reg__U594_in = delay_reg__U593_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U594 (
    .clk(delay_reg__U594_clk),
    .in(delay_reg__U594_in),
    .out(delay_reg__U594_out)
);
assign delay_reg__U595_clk = clk;
assign delay_reg__U595_in = delay_reg__U594_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U595 (
    .clk(delay_reg__U595_clk),
    .in(delay_reg__U595_in),
    .out(delay_reg__U595_out)
);
assign delay_reg__U596_clk = clk;
assign delay_reg__U596_in = delay_reg__U595_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U596 (
    .clk(delay_reg__U596_clk),
    .in(delay_reg__U596_in),
    .out(delay_reg__U596_out)
);
assign delay_reg__U597_clk = clk;
assign delay_reg__U597_in = delay_reg__U596_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U597 (
    .clk(delay_reg__U597_clk),
    .in(delay_reg__U597_in),
    .out(delay_reg__U597_out)
);
assign delay_reg__U598_clk = clk;
assign delay_reg__U598_in = delay_reg__U597_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U598 (
    .clk(delay_reg__U598_clk),
    .in(delay_reg__U598_in),
    .out(delay_reg__U598_out)
);
assign delay_reg__U599_clk = clk;
assign delay_reg__U599_in = delay_reg__U598_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U599 (
    .clk(delay_reg__U599_clk),
    .in(delay_reg__U599_in),
    .out(delay_reg__U599_out)
);
assign delay_reg__U600_clk = clk;
assign delay_reg__U600_in = delay_reg__U599_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U600 (
    .clk(delay_reg__U600_clk),
    .in(delay_reg__U600_in),
    .out(delay_reg__U600_out)
);
assign delay_reg__U601_clk = clk;
assign delay_reg__U601_in = delay_reg__U600_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U601 (
    .clk(delay_reg__U601_clk),
    .in(delay_reg__U601_in),
    .out(delay_reg__U601_out)
);
assign delay_reg__U602_clk = clk;
assign delay_reg__U602_in = delay_reg__U601_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U602 (
    .clk(delay_reg__U602_clk),
    .in(delay_reg__U602_in),
    .out(delay_reg__U602_out)
);
assign delay_reg__U603_clk = clk;
assign delay_reg__U603_in = delay_reg__U602_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U603 (
    .clk(delay_reg__U603_clk),
    .in(delay_reg__U603_in),
    .out(delay_reg__U603_out)
);
assign delay_reg__U604_clk = clk;
assign delay_reg__U604_in = delay_reg__U603_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U604 (
    .clk(delay_reg__U604_clk),
    .in(delay_reg__U604_in),
    .out(delay_reg__U604_out)
);
assign delay_reg__U605_clk = clk;
assign delay_reg__U605_in = delay_reg__U604_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U605 (
    .clk(delay_reg__U605_clk),
    .in(delay_reg__U605_in),
    .out(delay_reg__U605_out)
);
assign delay_reg__U95_clk = clk;
assign delay_reg__U95_in = op_hcompute_hw_output_stencil_port_controller_valid;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U95 (
    .clk(delay_reg__U95_clk),
    .in(delay_reg__U95_in),
    .out(delay_reg__U95_out)
);
assign delay_reg__U96_clk = clk;
assign delay_reg__U96_in = delay_reg__U95_out;
corebit_reg #(
    .clk_posedge(1'b1),
    .init(1'b0)
) delay_reg__U96 (
    .clk(delay_reg__U96_clk),
    .in(delay_reg__U96_in),
    .out(delay_reg__U96_out)
);
assign hw_input_global_wrapper_stencil_clk = clk;
assign hw_input_global_wrapper_stencil_flush = flush;
assign hw_input_global_wrapper_stencil_rst_n = rst_n;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen = op_hcompute_hw_input_global_wrapper_stencil_write_start_out;
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0] = op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write[0];
hw_input_global_wrapper_stencil_ub hw_input_global_wrapper_stencil (
    .clk(hw_input_global_wrapper_stencil_clk),
    .flush(hw_input_global_wrapper_stencil_flush),
    .rst_n(hw_input_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_input_global_wrapper_stencil_write_wen(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_input_global_wrapper_stencil_write(hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign hw_kernel_global_wrapper_stencil_clk = clk;
assign hw_kernel_global_wrapper_stencil_flush = flush;
assign hw_kernel_global_wrapper_stencil_rst_n = rst_n;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren = op_hcompute_conv_stencil_3_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren = op_hcompute_conv_stencil_4_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren = op_hcompute_conv_stencil_5_read_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out;
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[4] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[4];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[3] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[3];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[2] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[2];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[1] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[1];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars[0] = op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out[0];
assign hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0] = op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write[0];
hw_kernel_global_wrapper_stencil_ub hw_kernel_global_wrapper_stencil (
    .clk(hw_kernel_global_wrapper_stencil_clk),
    .flush(hw_kernel_global_wrapper_stencil_flush),
    .rst_n(hw_kernel_global_wrapper_stencil_rst_n),
    .op_hcompute_conv_stencil_3_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ren),
    .op_hcompute_conv_stencil_3_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read_ctrl_vars),
    .op_hcompute_conv_stencil_3_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .op_hcompute_conv_stencil_4_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ren),
    .op_hcompute_conv_stencil_4_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read_ctrl_vars),
    .op_hcompute_conv_stencil_4_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .op_hcompute_conv_stencil_5_read_ren(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ren),
    .op_hcompute_conv_stencil_5_read_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read_ctrl_vars),
    .op_hcompute_conv_stencil_5_read(hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_wen(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_wen),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write_ctrl_vars),
    .op_hcompute_hw_kernel_global_wrapper_stencil_write(hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_conv_stencil_clk = clk;
cu_op_hcompute_conv_stencil op_hcompute_conv_stencil (
    .clk(op_hcompute_conv_stencil_clk),
    .conv_stencil_op_hcompute_conv_stencil_write(op_hcompute_conv_stencil_conv_stencil_op_hcompute_conv_stencil_write)
);
assign op_hcompute_conv_stencil_1_clk = clk;
cu_op_hcompute_conv_stencil_1 op_hcompute_conv_stencil_1 (
    .clk(op_hcompute_conv_stencil_1_clk),
    .conv_stencil_op_hcompute_conv_stencil_1_write(op_hcompute_conv_stencil_1_conv_stencil_op_hcompute_conv_stencil_1_write)
);
assign op_hcompute_conv_stencil_1_exe_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_exe_start_pt__U42 op_hcompute_conv_stencil_1_exe_start (
    .in(op_hcompute_conv_stencil_1_exe_start_in),
    .out(op_hcompute_conv_stencil_1_exe_start_out)
);
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_exe_start_control_vars_pt__U43 op_hcompute_conv_stencil_1_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_1_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_port_controller_clk = clk;
affine_controller__U23 op_hcompute_conv_stencil_1_port_controller (
    .clk(op_hcompute_conv_stencil_1_port_controller_clk),
    .valid(op_hcompute_conv_stencil_1_port_controller_valid),
    .d(op_hcompute_conv_stencil_1_port_controller_d)
);
assign op_hcompute_conv_stencil_1_read_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_read_start_pt__U40 op_hcompute_conv_stencil_1_read_start (
    .in(op_hcompute_conv_stencil_1_read_start_in),
    .out(op_hcompute_conv_stencil_1_read_start_out)
);
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_read_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_read_start_control_vars_pt__U41 op_hcompute_conv_stencil_1_read_start_control_vars (
    .in(op_hcompute_conv_stencil_1_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_1_write_start_in = op_hcompute_conv_stencil_1_port_controller_valid;
op_hcompute_conv_stencil_1_write_start_pt__U44 op_hcompute_conv_stencil_1_write_start (
    .in(op_hcompute_conv_stencil_1_write_start_in),
    .out(op_hcompute_conv_stencil_1_write_start_out)
);
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[2] = op_hcompute_conv_stencil_1_port_controller_d[2];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[1] = op_hcompute_conv_stencil_1_port_controller_d[1];
assign op_hcompute_conv_stencil_1_write_start_control_vars_in[0] = op_hcompute_conv_stencil_1_port_controller_d[0];
op_hcompute_conv_stencil_1_write_start_control_vars_pt__U45 op_hcompute_conv_stencil_1_write_start_control_vars (
    .in(op_hcompute_conv_stencil_1_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_1_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_clk = clk;
cu_op_hcompute_conv_stencil_2 op_hcompute_conv_stencil_2 (
    .clk(op_hcompute_conv_stencil_2_clk),
    .conv_stencil_op_hcompute_conv_stencil_2_write(op_hcompute_conv_stencil_2_conv_stencil_op_hcompute_conv_stencil_2_write)
);
assign op_hcompute_conv_stencil_2_exe_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_exe_start_pt__U65 op_hcompute_conv_stencil_2_exe_start (
    .in(op_hcompute_conv_stencil_2_exe_start_in),
    .out(op_hcompute_conv_stencil_2_exe_start_out)
);
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_exe_start_control_vars_pt__U66 op_hcompute_conv_stencil_2_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_2_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_port_controller_clk = clk;
affine_controller__U46 op_hcompute_conv_stencil_2_port_controller (
    .clk(op_hcompute_conv_stencil_2_port_controller_clk),
    .valid(op_hcompute_conv_stencil_2_port_controller_valid),
    .d(op_hcompute_conv_stencil_2_port_controller_d)
);
assign op_hcompute_conv_stencil_2_read_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_read_start_pt__U63 op_hcompute_conv_stencil_2_read_start (
    .in(op_hcompute_conv_stencil_2_read_start_in),
    .out(op_hcompute_conv_stencil_2_read_start_out)
);
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_read_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_read_start_control_vars_pt__U64 op_hcompute_conv_stencil_2_read_start_control_vars (
    .in(op_hcompute_conv_stencil_2_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_2_write_start_in = op_hcompute_conv_stencil_2_port_controller_valid;
op_hcompute_conv_stencil_2_write_start_pt__U67 op_hcompute_conv_stencil_2_write_start (
    .in(op_hcompute_conv_stencil_2_write_start_in),
    .out(op_hcompute_conv_stencil_2_write_start_out)
);
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[2] = op_hcompute_conv_stencil_2_port_controller_d[2];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[1] = op_hcompute_conv_stencil_2_port_controller_d[1];
assign op_hcompute_conv_stencil_2_write_start_control_vars_in[0] = op_hcompute_conv_stencil_2_port_controller_d[0];
op_hcompute_conv_stencil_2_write_start_control_vars_pt__U68 op_hcompute_conv_stencil_2_write_start_control_vars (
    .in(op_hcompute_conv_stencil_2_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_2_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_clk = clk;
assign op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read[0] = conv_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[7];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[6];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[5];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[4];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[3];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[2];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[1];
assign op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read[0];
cu_op_hcompute_conv_stencil_3 op_hcompute_conv_stencil_3 (
    .clk(op_hcompute_conv_stencil_3_clk),
    .conv_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read(op_hcompute_conv_stencil_3_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_3_read),
    .conv_stencil_op_hcompute_conv_stencil_3_write(op_hcompute_conv_stencil_3_conv_stencil_op_hcompute_conv_stencil_3_write)
);
assign op_hcompute_conv_stencil_3_exe_start_in = delay_reg__U572_out;
op_hcompute_conv_stencil_3_exe_start_pt__U570 op_hcompute_conv_stencil_3_exe_start (
    .in(op_hcompute_conv_stencil_3_exe_start_in),
    .out(op_hcompute_conv_stencil_3_exe_start_out)
);
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[4] = arr__U581_out[4];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[3] = arr__U581_out[3];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[2] = arr__U581_out[2];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[1] = arr__U581_out[1];
assign op_hcompute_conv_stencil_3_exe_start_control_vars_in[0] = arr__U581_out[0];
op_hcompute_conv_stencil_3_exe_start_control_vars_pt__U573 op_hcompute_conv_stencil_3_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_3_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_port_controller_clk = clk;
affine_controller__U538 op_hcompute_conv_stencil_3_port_controller (
    .clk(op_hcompute_conv_stencil_3_port_controller_clk),
    .valid(op_hcompute_conv_stencil_3_port_controller_valid),
    .d(op_hcompute_conv_stencil_3_port_controller_d)
);
assign op_hcompute_conv_stencil_3_read_start_in = op_hcompute_conv_stencil_3_port_controller_valid;
op_hcompute_conv_stencil_3_read_start_pt__U568 op_hcompute_conv_stencil_3_read_start (
    .in(op_hcompute_conv_stencil_3_read_start_in),
    .out(op_hcompute_conv_stencil_3_read_start_out)
);
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[4] = op_hcompute_conv_stencil_3_port_controller_d[4];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[3] = op_hcompute_conv_stencil_3_port_controller_d[3];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[2] = op_hcompute_conv_stencil_3_port_controller_d[2];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[1] = op_hcompute_conv_stencil_3_port_controller_d[1];
assign op_hcompute_conv_stencil_3_read_start_control_vars_in[0] = op_hcompute_conv_stencil_3_port_controller_d[0];
op_hcompute_conv_stencil_3_read_start_control_vars_pt__U569 op_hcompute_conv_stencil_3_read_start_control_vars (
    .in(op_hcompute_conv_stencil_3_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_3_write_start_in = delay_reg__U605_out;
op_hcompute_conv_stencil_3_write_start_pt__U588 op_hcompute_conv_stencil_3_write_start (
    .in(op_hcompute_conv_stencil_3_write_start_in),
    .out(op_hcompute_conv_stencil_3_write_start_out)
);
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[4] = arr__U719_out[4];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[3] = arr__U719_out[3];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[2] = arr__U719_out[2];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[1] = arr__U719_out[1];
assign op_hcompute_conv_stencil_3_write_start_control_vars_in[0] = arr__U719_out[0];
op_hcompute_conv_stencil_3_write_start_control_vars_pt__U606 op_hcompute_conv_stencil_3_write_start_control_vars (
    .in(op_hcompute_conv_stencil_3_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_3_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_clk = clk;
assign op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read[0] = conv_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[7];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[6];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[5];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[4];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[3];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[2];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[1];
assign op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read[0];
cu_op_hcompute_conv_stencil_4 op_hcompute_conv_stencil_4 (
    .clk(op_hcompute_conv_stencil_4_clk),
    .conv_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read(op_hcompute_conv_stencil_4_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_4_read),
    .conv_stencil_op_hcompute_conv_stencil_4_write(op_hcompute_conv_stencil_4_conv_stencil_op_hcompute_conv_stencil_4_write)
);
assign op_hcompute_conv_stencil_4_exe_start_in = delay_reg__U384_out;
op_hcompute_conv_stencil_4_exe_start_pt__U382 op_hcompute_conv_stencil_4_exe_start (
    .in(op_hcompute_conv_stencil_4_exe_start_in),
    .out(op_hcompute_conv_stencil_4_exe_start_out)
);
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[4] = arr__U393_out[4];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[3] = arr__U393_out[3];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[2] = arr__U393_out[2];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[1] = arr__U393_out[1];
assign op_hcompute_conv_stencil_4_exe_start_control_vars_in[0] = arr__U393_out[0];
op_hcompute_conv_stencil_4_exe_start_control_vars_pt__U385 op_hcompute_conv_stencil_4_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_4_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_port_controller_clk = clk;
affine_controller__U350 op_hcompute_conv_stencil_4_port_controller (
    .clk(op_hcompute_conv_stencil_4_port_controller_clk),
    .valid(op_hcompute_conv_stencil_4_port_controller_valid),
    .d(op_hcompute_conv_stencil_4_port_controller_d)
);
assign op_hcompute_conv_stencil_4_read_start_in = op_hcompute_conv_stencil_4_port_controller_valid;
op_hcompute_conv_stencil_4_read_start_pt__U380 op_hcompute_conv_stencil_4_read_start (
    .in(op_hcompute_conv_stencil_4_read_start_in),
    .out(op_hcompute_conv_stencil_4_read_start_out)
);
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[4] = op_hcompute_conv_stencil_4_port_controller_d[4];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[3] = op_hcompute_conv_stencil_4_port_controller_d[3];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[2] = op_hcompute_conv_stencil_4_port_controller_d[2];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[1] = op_hcompute_conv_stencil_4_port_controller_d[1];
assign op_hcompute_conv_stencil_4_read_start_control_vars_in[0] = op_hcompute_conv_stencil_4_port_controller_d[0];
op_hcompute_conv_stencil_4_read_start_control_vars_pt__U381 op_hcompute_conv_stencil_4_read_start_control_vars (
    .in(op_hcompute_conv_stencil_4_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_4_write_start_in = delay_reg__U417_out;
op_hcompute_conv_stencil_4_write_start_pt__U400 op_hcompute_conv_stencil_4_write_start (
    .in(op_hcompute_conv_stencil_4_write_start_in),
    .out(op_hcompute_conv_stencil_4_write_start_out)
);
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[4] = arr__U531_out[4];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[3] = arr__U531_out[3];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[2] = arr__U531_out[2];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[1] = arr__U531_out[1];
assign op_hcompute_conv_stencil_4_write_start_control_vars_in[0] = arr__U531_out[0];
op_hcompute_conv_stencil_4_write_start_control_vars_pt__U418 op_hcompute_conv_stencil_4_write_start_control_vars (
    .in(op_hcompute_conv_stencil_4_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_4_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_clk = clk;
assign op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read[0] = conv_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[7];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[6];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[5];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[4];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[3];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[2];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[1];
assign op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0] = hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read[0];
cu_op_hcompute_conv_stencil_5 op_hcompute_conv_stencil_5 (
    .clk(op_hcompute_conv_stencil_5_clk),
    .conv_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_read),
    .hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_input_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read(op_hcompute_conv_stencil_5_hw_kernel_global_wrapper_stencil_op_hcompute_conv_stencil_5_read),
    .conv_stencil_op_hcompute_conv_stencil_5_write(op_hcompute_conv_stencil_5_conv_stencil_op_hcompute_conv_stencil_5_write)
);
assign op_hcompute_conv_stencil_5_exe_start_in = delay_reg__U160_out;
op_hcompute_conv_stencil_5_exe_start_pt__U158 op_hcompute_conv_stencil_5_exe_start (
    .in(op_hcompute_conv_stencil_5_exe_start_in),
    .out(op_hcompute_conv_stencil_5_exe_start_out)
);
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[4] = arr__U169_out[4];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[3] = arr__U169_out[3];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[2] = arr__U169_out[2];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[1] = arr__U169_out[1];
assign op_hcompute_conv_stencil_5_exe_start_control_vars_in[0] = arr__U169_out[0];
op_hcompute_conv_stencil_5_exe_start_control_vars_pt__U161 op_hcompute_conv_stencil_5_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_5_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_port_controller_clk = clk;
affine_controller__U126 op_hcompute_conv_stencil_5_port_controller (
    .clk(op_hcompute_conv_stencil_5_port_controller_clk),
    .valid(op_hcompute_conv_stencil_5_port_controller_valid),
    .d(op_hcompute_conv_stencil_5_port_controller_d)
);
assign op_hcompute_conv_stencil_5_read_start_in = op_hcompute_conv_stencil_5_port_controller_valid;
op_hcompute_conv_stencil_5_read_start_pt__U156 op_hcompute_conv_stencil_5_read_start (
    .in(op_hcompute_conv_stencil_5_read_start_in),
    .out(op_hcompute_conv_stencil_5_read_start_out)
);
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[4] = op_hcompute_conv_stencil_5_port_controller_d[4];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[3] = op_hcompute_conv_stencil_5_port_controller_d[3];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[2] = op_hcompute_conv_stencil_5_port_controller_d[2];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[1] = op_hcompute_conv_stencil_5_port_controller_d[1];
assign op_hcompute_conv_stencil_5_read_start_control_vars_in[0] = op_hcompute_conv_stencil_5_port_controller_d[0];
op_hcompute_conv_stencil_5_read_start_control_vars_pt__U157 op_hcompute_conv_stencil_5_read_start_control_vars (
    .in(op_hcompute_conv_stencil_5_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_5_write_start_in = delay_reg__U193_out;
op_hcompute_conv_stencil_5_write_start_pt__U176 op_hcompute_conv_stencil_5_write_start (
    .in(op_hcompute_conv_stencil_5_write_start_in),
    .out(op_hcompute_conv_stencil_5_write_start_out)
);
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[4] = arr__U307_out[4];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[3] = arr__U307_out[3];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[2] = arr__U307_out[2];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[1] = arr__U307_out[1];
assign op_hcompute_conv_stencil_5_write_start_control_vars_in[0] = arr__U307_out[0];
op_hcompute_conv_stencil_5_write_start_control_vars_pt__U194 op_hcompute_conv_stencil_5_write_start_control_vars (
    .in(op_hcompute_conv_stencil_5_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_5_write_start_control_vars_out)
);
assign op_hcompute_conv_stencil_exe_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_exe_start_pt__U19 op_hcompute_conv_stencil_exe_start (
    .in(op_hcompute_conv_stencil_exe_start_in),
    .out(op_hcompute_conv_stencil_exe_start_out)
);
assign op_hcompute_conv_stencil_exe_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_exe_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_exe_start_control_vars_pt__U20 op_hcompute_conv_stencil_exe_start_control_vars (
    .in(op_hcompute_conv_stencil_exe_start_control_vars_in),
    .out(op_hcompute_conv_stencil_exe_start_control_vars_out)
);
assign op_hcompute_conv_stencil_port_controller_clk = clk;
affine_controller__U0 op_hcompute_conv_stencil_port_controller (
    .clk(op_hcompute_conv_stencil_port_controller_clk),
    .valid(op_hcompute_conv_stencil_port_controller_valid),
    .d(op_hcompute_conv_stencil_port_controller_d)
);
assign op_hcompute_conv_stencil_read_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_read_start_pt__U17 op_hcompute_conv_stencil_read_start (
    .in(op_hcompute_conv_stencil_read_start_in),
    .out(op_hcompute_conv_stencil_read_start_out)
);
assign op_hcompute_conv_stencil_read_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_read_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_read_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_read_start_control_vars_pt__U18 op_hcompute_conv_stencil_read_start_control_vars (
    .in(op_hcompute_conv_stencil_read_start_control_vars_in),
    .out(op_hcompute_conv_stencil_read_start_control_vars_out)
);
assign op_hcompute_conv_stencil_write_start_in = op_hcompute_conv_stencil_port_controller_valid;
op_hcompute_conv_stencil_write_start_pt__U21 op_hcompute_conv_stencil_write_start (
    .in(op_hcompute_conv_stencil_write_start_in),
    .out(op_hcompute_conv_stencil_write_start_out)
);
assign op_hcompute_conv_stencil_write_start_control_vars_in[2] = op_hcompute_conv_stencil_port_controller_d[2];
assign op_hcompute_conv_stencil_write_start_control_vars_in[1] = op_hcompute_conv_stencil_port_controller_d[1];
assign op_hcompute_conv_stencil_write_start_control_vars_in[0] = op_hcompute_conv_stencil_port_controller_d[0];
op_hcompute_conv_stencil_write_start_control_vars_pt__U22 op_hcompute_conv_stencil_write_start_control_vars (
    .in(op_hcompute_conv_stencil_write_start_control_vars_in),
    .out(op_hcompute_conv_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0] = hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_input_global_wrapper_stencil op_hcompute_hw_input_global_wrapper_stencil (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_clk),
    .hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read(op_hcompute_hw_input_global_wrapper_stencil_hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read),
    .hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write(op_hcompute_hw_input_global_wrapper_stencil_hw_input_global_wrapper_stencil_op_hcompute_hw_input_global_wrapper_stencil_write)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_exe_start_pt__U751 op_hcompute_hw_input_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_pt__U752 op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U726 op_hcompute_hw_input_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_input_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_input_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_read_start_pt__U749 op_hcompute_hw_input_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_in),
    .out(hw_input_stencil_op_hcompute_hw_input_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_pt__U750 op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_in = op_hcompute_hw_input_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_input_global_wrapper_stencil_write_start_pt__U753 op_hcompute_hw_input_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_input_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_pt__U754 op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_input_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_clk = clk;
assign op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0] = hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read[0];
cu_op_hcompute_hw_kernel_global_wrapper_stencil op_hcompute_hw_kernel_global_wrapper_stencil (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_clk),
    .hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read),
    .hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write(op_hcompute_hw_kernel_global_wrapper_stencil_hw_kernel_global_wrapper_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_write)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_pt__U346 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_pt__U347 op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk = clk;
affine_controller__U314 op_hcompute_hw_kernel_global_wrapper_stencil_port_controller (
    .clk(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_clk),
    .valid(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid),
    .d(op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_pt__U344 op_hcompute_hw_kernel_global_wrapper_stencil_read_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_in),
    .out(hw_kernel_stencil_op_hcompute_hw_kernel_global_wrapper_stencil_read_en)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_pt__U345 op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_valid;
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_pt__U348 op_hcompute_hw_kernel_global_wrapper_stencil_write_start (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_out)
);
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[4] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[4];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[3] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[3];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[2] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[2];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[1] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[1];
assign op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in[0] = op_hcompute_hw_kernel_global_wrapper_stencil_port_controller_d[0];
op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_pt__U349 op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars (
    .in(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_kernel_global_wrapper_stencil_write_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_clk = clk;
assign op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read[0] = conv_stencil_op_hcompute_hw_output_stencil_read[0];
cu_op_hcompute_hw_output_stencil op_hcompute_hw_output_stencil (
    .clk(op_hcompute_hw_output_stencil_clk),
    .conv_stencil_op_hcompute_hw_output_stencil_read(op_hcompute_hw_output_stencil_conv_stencil_op_hcompute_hw_output_stencil_read),
    .hw_output_stencil_op_hcompute_hw_output_stencil_write(op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write)
);
assign op_hcompute_hw_output_stencil_exe_start_in = delay_reg__U96_out;
op_hcompute_hw_output_stencil_exe_start_pt__U94 op_hcompute_hw_output_stencil_exe_start (
    .in(op_hcompute_hw_output_stencil_exe_start_in),
    .out(op_hcompute_hw_output_stencil_exe_start_out)
);
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[3] = arr__U104_out[3];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[2] = arr__U104_out[2];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[1] = arr__U104_out[1];
assign op_hcompute_hw_output_stencil_exe_start_control_vars_in[0] = arr__U104_out[0];
op_hcompute_hw_output_stencil_exe_start_control_vars_pt__U97 op_hcompute_hw_output_stencil_exe_start_control_vars (
    .in(op_hcompute_hw_output_stencil_exe_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_exe_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_port_controller_clk = clk;
affine_controller__U69 op_hcompute_hw_output_stencil_port_controller (
    .clk(op_hcompute_hw_output_stencil_port_controller_clk),
    .valid(op_hcompute_hw_output_stencil_port_controller_valid),
    .d(op_hcompute_hw_output_stencil_port_controller_d)
);
assign op_hcompute_hw_output_stencil_read_start_in = op_hcompute_hw_output_stencil_port_controller_valid;
op_hcompute_hw_output_stencil_read_start_pt__U92 op_hcompute_hw_output_stencil_read_start (
    .in(op_hcompute_hw_output_stencil_read_start_in),
    .out(op_hcompute_hw_output_stencil_read_start_out)
);
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[3] = op_hcompute_hw_output_stencil_port_controller_d[3];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[2] = op_hcompute_hw_output_stencil_port_controller_d[2];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[1] = op_hcompute_hw_output_stencil_port_controller_d[1];
assign op_hcompute_hw_output_stencil_read_start_control_vars_in[0] = op_hcompute_hw_output_stencil_port_controller_d[0];
op_hcompute_hw_output_stencil_read_start_control_vars_pt__U93 op_hcompute_hw_output_stencil_read_start_control_vars (
    .in(op_hcompute_hw_output_stencil_read_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_read_start_control_vars_out)
);
assign op_hcompute_hw_output_stencil_write_start_in = delay_reg__U112_out;
op_hcompute_hw_output_stencil_write_start_pt__U110 op_hcompute_hw_output_stencil_write_start (
    .in(op_hcompute_hw_output_stencil_write_start_in),
    .out(hw_output_stencil_op_hcompute_hw_output_stencil_write_valid)
);
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[3] = arr__U120_out[3];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[2] = arr__U120_out[2];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[1] = arr__U120_out[1];
assign op_hcompute_hw_output_stencil_write_start_control_vars_in[0] = arr__U120_out[0];
op_hcompute_hw_output_stencil_write_start_control_vars_pt__U113 op_hcompute_hw_output_stencil_write_start_control_vars (
    .in(op_hcompute_hw_output_stencil_write_start_control_vars_in),
    .out(op_hcompute_hw_output_stencil_write_start_control_vars_out)
);
assign hw_output_stencil_op_hcompute_hw_output_stencil_write[0] = op_hcompute_hw_output_stencil_hw_output_stencil_op_hcompute_hw_output_stencil_write[0];
endmodule

